module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_017_not;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_063_not;
  wire cgp_core_064;
  wire cgp_core_065;

  assign cgp_core_014 = ~(input_e[1] ^ input_d[0]);
  assign cgp_core_016 = input_a[1] | input_a[1];
  assign cgp_core_017_not = ~input_f[0];
  assign cgp_core_019 = input_c[1] ^ input_c[0];
  assign cgp_core_021 = input_c[0] ^ input_b[0];
  assign cgp_core_022 = ~(input_d[1] & input_e[1]);
  assign cgp_core_024 = input_e[0] & input_f[0];
  assign cgp_core_025 = input_e[0] ^ input_c[0];
  assign cgp_core_026 = ~input_e[1];
  assign cgp_core_027 = ~input_c[0];
  assign cgp_core_029 = ~(input_c[1] | input_f[1]);
  assign cgp_core_032 = ~(input_d[0] | cgp_core_029);
  assign cgp_core_033 = ~(input_e[1] ^ input_f[1]);
  assign cgp_core_035 = ~(input_b[1] | input_e[0]);
  assign cgp_core_036 = input_b[0] ^ input_a[1];
  assign cgp_core_037 = ~input_e[0];
  assign cgp_core_038 = cgp_core_025 ^ input_c[1];
  assign cgp_core_039 = input_f[0] ^ input_f[0];
  assign cgp_core_040 = input_c[0] & input_a[1];
  assign cgp_core_041 = input_d[0] | cgp_core_040;
  assign cgp_core_042 = input_d[0] | input_f[0];
  assign cgp_core_044 = input_a[1] ^ input_e[1];
  assign cgp_core_045 = input_c[0] ^ input_c[0];
  assign cgp_core_046 = input_c[1] & input_a[0];
  assign cgp_core_048 = input_c[0] ^ input_a[0];
  assign cgp_core_050 = input_d[1] ^ input_b[1];
  assign cgp_core_052 = ~(input_d[0] ^ input_a[1]);
  assign cgp_core_053_not = ~input_d[1];
  assign cgp_core_054 = ~input_a[1];
  assign cgp_core_055 = ~(input_d[1] & input_d[1]);
  assign cgp_core_058 = ~(input_c[1] & input_f[0]);
  assign cgp_core_059 = input_b[1] & input_c[0];
  assign cgp_core_063_not = ~input_d[1];
  assign cgp_core_064 = ~(input_f[0] | input_e[0]);
  assign cgp_core_065 = ~(input_b[1] & input_d[1]);

  assign cgp_out[0] = 1'b0;
endmodule