module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_037_not;
  wire cgp_core_039_not;
  wire cgp_core_043;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_016 = input_a[0] ^ input_d[1];
  assign cgp_core_017 = input_a[0] & input_c[0];
  assign cgp_core_018 = input_a[1] ^ input_c[1];
  assign cgp_core_019 = input_a[1] & input_c[1];
  assign cgp_core_020 = cgp_core_018 ^ input_g[1];
  assign cgp_core_021 = cgp_core_018 & input_d[0];
  assign cgp_core_023 = input_e[0] ^ input_g[0];
  assign cgp_core_024 = input_e[0] & input_g[0];
  assign cgp_core_025 = input_g[0] ^ input_g[1];
  assign cgp_core_026 = input_e[1] & input_d[0];
  assign cgp_core_027 = cgp_core_025 ^ input_g[0];
  assign cgp_core_031 = input_d[0] & cgp_core_023;
  assign cgp_core_032 = input_d[1] | cgp_core_027;
  assign cgp_core_034 = cgp_core_032 ^ input_b[0];
  assign cgp_core_037_not = ~cgp_core_026;
  assign cgp_core_039_not = ~cgp_core_016;
  assign cgp_core_043 = cgp_core_020 ^ cgp_core_016;
  assign cgp_core_053 = input_b[0] ^ input_f[0];
  assign cgp_core_054 = input_b[0] & input_b[0];
  assign cgp_core_055 = input_b[1] ^ input_f[1];
  assign cgp_core_056 = input_b[1] & input_f[1];
  assign cgp_core_063 = input_f[1] & input_c[0];
  assign cgp_core_064 = cgp_core_056 ^ cgp_core_056;
  assign cgp_core_067 = ~(input_b[0] ^ input_a[1]);
  assign cgp_core_073 = input_a[0] & input_d[0];
  assign cgp_core_074 = ~input_c[0];
  assign cgp_core_075 = cgp_core_039_not & cgp_core_074;
  assign cgp_core_077 = ~(cgp_core_039_not ^ cgp_core_053);
  assign cgp_core_078 = input_b[1] & cgp_core_073;

  assign cgp_out[0] = 1'b1;
endmodule