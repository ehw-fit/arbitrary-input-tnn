module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_108;
  wire cgp_core_109;

  assign cgp_core_020 = ~input_g[0];
  assign cgp_core_021 = input_c[1] & input_i[0];
  assign cgp_core_022 = input_i[1] | input_h[1];
  assign cgp_core_023 = input_h[1] & input_i[1];
  assign cgp_core_027 = ~input_h[1];
  assign cgp_core_028 = ~input_g[1];
  assign cgp_core_029 = ~(input_b[0] | input_b[0]);
  assign cgp_core_030 = input_d[1] & cgp_core_022;
  assign cgp_core_031 = input_h[0] ^ input_c[1];
  assign cgp_core_032 = ~input_e[1];
  assign cgp_core_034 = cgp_core_023 | cgp_core_030;
  assign cgp_core_035 = input_a[1] ^ input_a[1];
  assign cgp_core_037 = input_i[1] & input_h[0];
  assign cgp_core_038 = input_b[1] & input_h[0];
  assign cgp_core_040 = input_g[1] ^ input_a[0];
  assign cgp_core_041 = input_c[1] & input_a[1];
  assign cgp_core_042 = input_g[1] | cgp_core_041;
  assign cgp_core_043 = ~input_e[0];
  assign cgp_core_044 = input_f[0] & input_d[1];
  assign cgp_core_047 = input_a[0] | input_a[0];
  assign cgp_core_049 = ~(input_a[1] | input_b[0]);
  assign cgp_core_050 = input_e[0] | input_b[0];
  assign cgp_core_052 = input_a[0] ^ input_g[0];
  assign cgp_core_054 = ~(input_h[0] | input_b[0]);
  assign cgp_core_055 = input_a[0] ^ input_d[0];
  assign cgp_core_056 = input_h[1] ^ input_d[0];
  assign cgp_core_057 = input_d[1] | input_i[0];
  assign cgp_core_059 = input_f[1] ^ input_i[0];
  assign cgp_core_062 = input_c[1] ^ input_c[1];
  assign cgp_core_067 = input_c[1] ^ input_f[0];
  assign cgp_core_068 = input_g[0] & input_a[1];
  assign cgp_core_069 = ~(input_f[0] & input_f[0]);
  assign cgp_core_070 = ~(input_e[1] ^ input_g[0]);
  assign cgp_core_071 = ~(input_e[0] & input_b[0]);
  assign cgp_core_072 = ~(input_a[0] | input_f[0]);
  assign cgp_core_073 = input_c[1] ^ input_e[1];
  assign cgp_core_074 = ~(input_e[0] & input_c[1]);
  assign cgp_core_076 = cgp_core_050 & input_f[1];
  assign cgp_core_080 = cgp_core_042 | input_e[1];
  assign cgp_core_081 = ~input_i[0];
  assign cgp_core_082 = cgp_core_080 | cgp_core_076;
  assign cgp_core_085 = input_d[0] & input_h[1];
  assign cgp_core_086 = input_h[1] | input_f[0];
  assign cgp_core_087 = ~input_e[1];
  assign cgp_core_088 = ~input_i[0];
  assign cgp_core_090 = ~(input_b[1] | cgp_core_082);
  assign cgp_core_092 = ~(input_d[1] ^ input_f[0]);
  assign cgp_core_094 = cgp_core_034 & cgp_core_090;
  assign cgp_core_095 = ~input_e[0];
  assign cgp_core_096 = input_c[0] ^ input_f[1];
  assign cgp_core_098 = input_d[1] & input_b[0];
  assign cgp_core_099 = ~(input_c[0] | input_h[0]);
  assign cgp_core_100 = input_a[0] ^ input_g[1];
  assign cgp_core_104 = ~input_a[1];
  assign cgp_core_105 = ~(input_d[1] & input_d[0]);
  assign cgp_core_106 = ~(input_g[0] | input_a[0]);
  assign cgp_core_107 = ~(input_i[0] | input_d[1]);
  assign cgp_core_108 = ~(input_h[1] ^ input_a[0]);
  assign cgp_core_109 = input_i[1] & input_c[0];

  assign cgp_out[0] = cgp_core_094;
endmodule