module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_015 = input_c[2] ^ input_d[0];
  assign cgp_core_016 = ~input_b[2];
  assign cgp_core_019 = ~input_c[0];
  assign cgp_core_020 = input_a[1] | input_b[1];
  assign cgp_core_021 = input_a[2] ^ input_b[2];
  assign cgp_core_022 = input_a[2] & input_b[2];
  assign cgp_core_023 = cgp_core_021 ^ cgp_core_020;
  assign cgp_core_024 = cgp_core_021 & cgp_core_020;
  assign cgp_core_025 = cgp_core_022 | cgp_core_024;
  assign cgp_core_026 = input_d[2] & input_b[0];
  assign cgp_core_027 = ~input_d[0];
  assign cgp_core_028 = ~(input_d[2] & input_b[0]);
  assign cgp_core_029 = input_c[1] & input_d[1];
  assign cgp_core_030 = input_c[0] & input_d[0];
  assign cgp_core_033 = input_c[2] ^ input_d[2];
  assign cgp_core_034 = input_c[2] & input_d[2];
  assign cgp_core_035 = cgp_core_033 ^ cgp_core_029;
  assign cgp_core_036 = cgp_core_033 & cgp_core_029;
  assign cgp_core_037 = cgp_core_034 | cgp_core_036;
  assign cgp_core_038 = ~cgp_core_037;
  assign cgp_core_039 = cgp_core_025 & cgp_core_038;
  assign cgp_core_040 = ~(cgp_core_025 ^ cgp_core_037);
  assign cgp_core_041 = ~cgp_core_035;
  assign cgp_core_042 = cgp_core_023 & cgp_core_041;
  assign cgp_core_043 = cgp_core_042 & cgp_core_040;
  assign cgp_core_045 = ~input_d[2];
  assign cgp_core_046 = input_a[1] | input_c[0];
  assign cgp_core_048 = ~(input_c[1] ^ input_d[0]);
  assign cgp_core_050_not = ~input_c[2];
  assign cgp_core_051 = ~(input_b[0] ^ input_b[0]);
  assign cgp_core_052 = ~(input_b[1] ^ input_d[1]);
  assign cgp_core_053_not = ~input_b[1];
  assign cgp_core_054 = ~input_c[2];
  assign cgp_core_058 = cgp_core_043 | cgp_core_039;
  assign cgp_core_059 = ~(input_c[0] ^ input_d[2]);

  assign cgp_out[0] = cgp_core_058;
endmodule