module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065_not;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_080;

  assign cgp_core_018 = input_a[0] & input_b[0];
  assign cgp_core_019 = input_a[1] | input_b[1];
  assign cgp_core_020 = input_a[1] & input_b[1];
  assign cgp_core_021 = ~(input_e[0] | input_e[2]);
  assign cgp_core_022 = cgp_core_019 & cgp_core_018;
  assign cgp_core_023 = cgp_core_020 | cgp_core_022;
  assign cgp_core_024 = input_a[2] ^ input_b[2];
  assign cgp_core_025 = input_a[2] & input_b[2];
  assign cgp_core_026 = cgp_core_024 ^ cgp_core_023;
  assign cgp_core_027 = cgp_core_024 & cgp_core_023;
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_032 = input_d[1] & input_c[1];
  assign cgp_core_036 = input_d[2] ^ input_e[2];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038 = cgp_core_036 ^ cgp_core_032;
  assign cgp_core_039 = cgp_core_036 & cgp_core_032;
  assign cgp_core_040 = cgp_core_037 | cgp_core_039;
  assign cgp_core_044 = input_a[1] ^ input_d[0];
  assign cgp_core_047 = ~input_d[0];
  assign cgp_core_048 = input_c[2] ^ cgp_core_038;
  assign cgp_core_050 = ~cgp_core_048;
  assign cgp_core_052 = input_c[2] | cgp_core_048;
  assign cgp_core_053 = cgp_core_040 | cgp_core_052;
  assign cgp_core_054 = cgp_core_040 & cgp_core_052;
  assign cgp_core_055 = input_a[1] ^ input_b[0];
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_057 = ~cgp_core_053;
  assign cgp_core_058 = cgp_core_028 & cgp_core_057;
  assign cgp_core_060 = ~(cgp_core_028 ^ cgp_core_053);
  assign cgp_core_061 = cgp_core_060 & cgp_core_056;
  assign cgp_core_062 = ~input_d[0];
  assign cgp_core_064 = cgp_core_026 & cgp_core_061;
  assign cgp_core_065_not = ~cgp_core_050;
  assign cgp_core_066 = cgp_core_065_not & cgp_core_061;
  assign cgp_core_067 = input_a[0] & input_b[2];
  assign cgp_core_068 = input_c[0] ^ input_c[2];
  assign cgp_core_070 = ~(input_e[0] & input_b[0]);
  assign cgp_core_073 = input_e[1] | input_c[2];
  assign cgp_core_074 = ~input_c[1];
  assign cgp_core_076 = ~(input_a[0] | input_c[0]);
  assign cgp_core_077 = cgp_core_066 | cgp_core_064;
  assign cgp_core_080 = cgp_core_077 | cgp_core_058;

  assign cgp_out[0] = cgp_core_080;
endmodule