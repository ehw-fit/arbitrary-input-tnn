module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030_not;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_078;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_086;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_096;
  wire cgp_core_097;

  assign cgp_core_018 = input_h[1] | input_c[0];
  assign cgp_core_019 = ~(input_f[1] & input_a[1]);
  assign cgp_core_020 = input_b[1] | input_c[1];
  assign cgp_core_021 = input_b[1] & input_c[1];
  assign cgp_core_025 = ~(input_c[0] | input_a[0]);
  assign cgp_core_026 = ~(input_e[1] ^ input_e[0]);
  assign cgp_core_028 = input_a[1] & cgp_core_020;
  assign cgp_core_029 = ~(input_h[0] | input_c[0]);
  assign cgp_core_030_not = ~input_h[0];
  assign cgp_core_032 = cgp_core_021 | cgp_core_028;
  assign cgp_core_034 = input_c[0] ^ input_b[1];
  assign cgp_core_035 = input_c[0] & input_g[0];
  assign cgp_core_036 = input_g[1] | input_h[1];
  assign cgp_core_037 = ~(input_c[1] ^ input_a[1]);
  assign cgp_core_038 = cgp_core_036 | cgp_core_035;
  assign cgp_core_039 = cgp_core_036 & input_g[0];
  assign cgp_core_041 = input_c[1] | input_f[0];
  assign cgp_core_043 = input_d[1] | cgp_core_038;
  assign cgp_core_044 = input_d[1] & cgp_core_038;
  assign cgp_core_045 = ~input_f[1];
  assign cgp_core_046 = cgp_core_043 & input_d[0];
  assign cgp_core_047 = cgp_core_044 | cgp_core_046;
  assign cgp_core_048 = cgp_core_039 | cgp_core_047;
  assign cgp_core_049 = input_h[1] & input_g[1];
  assign cgp_core_050 = input_f[1] | input_a[0];
  assign cgp_core_052 = ~input_h[1];
  assign cgp_core_054 = ~input_b[0];
  assign cgp_core_055 = input_d[0] | input_h[1];
  assign cgp_core_059 = ~(input_e[1] & input_b[1]);
  assign cgp_core_061 = cgp_core_048 | cgp_core_032;
  assign cgp_core_064 = cgp_core_049 | cgp_core_061;
  assign cgp_core_065 = input_d[1] & input_d[1];
  assign cgp_core_067 = input_c[1] | input_a[1];
  assign cgp_core_068 = input_e[0] & input_f[0];
  assign cgp_core_069 = input_e[1] ^ input_f[1];
  assign cgp_core_070 = input_e[1] & input_f[1];
  assign cgp_core_071 = cgp_core_069 ^ input_f[0];
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~(input_c[1] | input_h[1]);
  assign cgp_core_078 = ~cgp_core_073;
  assign cgp_core_081 = input_a[0] & input_d[1];
  assign cgp_core_082 = input_e[0] & input_c[0];
  assign cgp_core_083 = ~(input_h[1] & input_d[1]);
  assign cgp_core_086 = ~(cgp_core_054 | cgp_core_071);
  assign cgp_core_089 = ~(input_e[1] & input_b[1]);
  assign cgp_core_090 = ~(input_d[1] | input_f[0]);
  assign cgp_core_092 = input_h[0] & cgp_core_086;
  assign cgp_core_096 = cgp_core_064 | cgp_core_092;
  assign cgp_core_097 = cgp_core_078 | cgp_core_096;

  assign cgp_out[0] = cgp_core_097;
endmodule