module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;

  assign cgp_core_020 = input_a[0] ^ input_b[0];
  assign cgp_core_021 = input_e[2] & input_b[0];
  assign cgp_core_023 = input_a[1] & input_b[1];
  assign cgp_core_024 = input_f[0] ^ input_a[0];
  assign cgp_core_027 = input_a[2] ^ input_b[2];
  assign cgp_core_028 = input_a[2] & input_b[2];
  assign cgp_core_029 = cgp_core_027 ^ input_f[2];
  assign cgp_core_031 = cgp_core_028 | input_b[1];
  assign cgp_core_032 = input_b[1] ^ input_d[0];
  assign cgp_core_033 = input_c[0] & input_d[0];
  assign cgp_core_034 = input_c[1] ^ input_d[1];
  assign cgp_core_035 = input_c[0] & input_d[1];
  assign cgp_core_036 = input_f[2] ^ input_c[0];
  assign cgp_core_037 = input_b[1] & input_b[1];
  assign cgp_core_038 = cgp_core_035 | cgp_core_037;
  assign cgp_core_039 = input_b[1] ^ input_d[2];
  assign cgp_core_041 = cgp_core_039 ^ cgp_core_038;
  assign cgp_core_042 = input_f[1] & cgp_core_038;
  assign cgp_core_043 = input_c[2] | cgp_core_042;
  assign cgp_core_044 = input_c[0] ^ input_f[0];
  assign cgp_core_045 = input_a[0] & input_c[0];
  assign cgp_core_046 = input_e[1] ^ input_f[1];
  assign cgp_core_047 = input_e[1] & input_f[1];
  assign cgp_core_048 = ~cgp_core_046;
  assign cgp_core_049 = cgp_core_046 & cgp_core_045;
  assign cgp_core_050 = cgp_core_047 | cgp_core_049;
  assign cgp_core_051 = input_c[1] ^ input_f[2];
  assign cgp_core_052 = input_e[2] & input_a[0];
  assign cgp_core_053 = cgp_core_051 ^ cgp_core_050;
  assign cgp_core_054 = input_a[2] & cgp_core_050;
  assign cgp_core_055 = cgp_core_052 | input_c[0];
  assign cgp_core_056 = ~cgp_core_032;
  assign cgp_core_057 = cgp_core_032 & cgp_core_044;
  assign cgp_core_058 = ~(cgp_core_036 & cgp_core_048);
  assign cgp_core_059 = cgp_core_036 & cgp_core_048;
  assign cgp_core_060 = cgp_core_058 ^ cgp_core_057;
  assign cgp_core_061 = cgp_core_058 & cgp_core_057;
  assign cgp_core_062 = cgp_core_059 | input_e[0];
  assign cgp_core_063 = cgp_core_041 ^ input_d[2];
  assign cgp_core_064 = cgp_core_041 & input_f[0];
  assign cgp_core_065 = input_d[0] ^ cgp_core_062;
  assign cgp_core_069 = cgp_core_043 & input_e[0];
  assign cgp_core_070 = ~input_f[2];
  assign cgp_core_071 = input_f[2] & cgp_core_064;
  assign cgp_core_072 = input_e[0] | cgp_core_071;
  assign cgp_core_073 = ~input_b[2];
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_078 = ~(cgp_core_031 ^ input_f[0]);
  assign cgp_core_080 = ~input_e[0];
  assign cgp_core_081 = cgp_core_029 & cgp_core_080;
  assign cgp_core_083 = ~(input_f[0] ^ input_c[2]);
  assign cgp_core_085 = ~input_f[0];
  assign cgp_core_086 = input_c[0] & input_f[2];
  assign cgp_core_090 = ~cgp_core_056;
  assign cgp_core_091 = cgp_core_020 & cgp_core_090;
  assign cgp_core_093 = ~(cgp_core_020 ^ cgp_core_056);

  assign cgp_out[0] = 1'b0;
endmodule