module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_015_not;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_026_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030_not;
  wire cgp_core_031_not;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_053;

  assign cgp_core_012 = ~(input_a[0] & input_d[1]);
  assign cgp_core_015_not = ~input_d[1];
  assign cgp_core_016 = ~(input_e[1] & input_a[1]);
  assign cgp_core_017 = input_d[1] ^ input_c[1];
  assign cgp_core_020 = ~input_e[0];
  assign cgp_core_021 = input_c[1] & input_c[0];
  assign cgp_core_026_not = ~input_d[1];
  assign cgp_core_028 = input_b[1] & input_d[0];
  assign cgp_core_029 = input_e[0] | input_c[0];
  assign cgp_core_030_not = ~input_a[1];
  assign cgp_core_031_not = ~input_e[0];
  assign cgp_core_034 = ~(input_c[1] | input_d[1]);
  assign cgp_core_035 = ~(input_e[1] | input_c[1]);
  assign cgp_core_037 = ~input_e[0];
  assign cgp_core_038 = input_a[1] & input_d[1];
  assign cgp_core_040 = input_d[0] ^ input_c[1];
  assign cgp_core_042 = ~(input_c[1] | input_e[0]);
  assign cgp_core_044 = ~input_a[0];
  assign cgp_core_045 = ~input_d[0];
  assign cgp_core_047 = ~input_b[1];
  assign cgp_core_050 = input_c[0] ^ input_d[0];
  assign cgp_core_053 = input_a[0] | input_d[0];

  assign cgp_out[0] = cgp_core_035;
endmodule