module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_022_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_081;
  wire cgp_core_086;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_095;
  wire cgp_core_096;

  assign cgp_core_020 = input_e[1] & input_c[0];
  assign cgp_core_022_not = ~input_f[0];
  assign cgp_core_024 = ~(input_g[1] ^ input_c[0]);
  assign cgp_core_025 = ~(input_b[0] ^ input_c[0]);
  assign cgp_core_026_not = ~input_b[1];
  assign cgp_core_028 = ~(input_d[1] & input_b[1]);
  assign cgp_core_029 = ~(input_f[0] & input_h[1]);
  assign cgp_core_030 = input_c[0] ^ input_a[1];
  assign cgp_core_031 = input_c[0] | input_h[0];
  assign cgp_core_032 = input_g[1] & input_d[1];
  assign cgp_core_033 = input_a[1] & input_h[1];
  assign cgp_core_034 = ~(input_h[0] ^ input_d[0]);
  assign cgp_core_037 = ~(input_f[1] & input_a[1]);
  assign cgp_core_040 = ~(input_b[0] ^ input_b[1]);
  assign cgp_core_041 = ~(input_f[0] | input_f[0]);
  assign cgp_core_043 = input_f[1] | input_g[1];
  assign cgp_core_044 = input_f[1] & input_g[1];
  assign cgp_core_046 = cgp_core_043 & input_b[1];
  assign cgp_core_047 = cgp_core_044 | cgp_core_046;
  assign cgp_core_048 = input_e[0] | input_f[0];
  assign cgp_core_050 = ~(input_c[0] ^ input_f[1]);
  assign cgp_core_051 = input_e[1] & input_c[1];
  assign cgp_core_052 = ~(input_f[1] ^ input_b[0]);
  assign cgp_core_053 = input_b[1] | input_a[1];
  assign cgp_core_055 = cgp_core_047 | cgp_core_051;
  assign cgp_core_057 = ~(input_h[0] ^ input_a[1]);
  assign cgp_core_059 = ~input_d[1];
  assign cgp_core_060 = input_a[0] | input_h[0];
  assign cgp_core_062 = input_d[1] ^ input_e[0];
  assign cgp_core_063 = ~(input_b[0] | input_f[0]);
  assign cgp_core_065 = input_a[1] & input_a[0];
  assign cgp_core_070 = input_c[0] | input_b[1];
  assign cgp_core_071 = input_f[0] & input_g[1];
  assign cgp_core_073 = ~cgp_core_055;
  assign cgp_core_074 = cgp_core_033 & cgp_core_073;
  assign cgp_core_075 = input_a[1] ^ input_d[1];
  assign cgp_core_077 = ~(input_b[0] & input_c[1]);
  assign cgp_core_081 = input_g[1] | input_f[1];
  assign cgp_core_086 = input_d[0] | input_b[1];
  assign cgp_core_089 = input_f[1] & input_e[1];
  assign cgp_core_090 = ~(input_f[1] ^ input_h[0]);
  assign cgp_core_092 = ~(input_e[0] ^ input_d[1]);
  assign cgp_core_095 = input_d[0] | input_g[0];
  assign cgp_core_096 = ~(input_h[0] & input_b[1]);

  assign cgp_out[0] = cgp_core_074;
endmodule