module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017 = ~input_e[0];
  assign cgp_core_018 = ~(input_d[0] & input_b[0]);
  assign cgp_core_019 = ~input_b[2];
  assign cgp_core_022 = input_c[1] & input_e[1];
  assign cgp_core_023 = input_c[2] | cgp_core_022;
  assign cgp_core_024 = ~(input_c[2] | input_e[1]);
  assign cgp_core_025 = input_c[2] & input_e[2];
  assign cgp_core_026 = input_e[2] | cgp_core_023;
  assign cgp_core_027_not = ~input_c[2];
  assign cgp_core_030 = ~(input_e[2] & input_c[0]);
  assign cgp_core_031 = ~(input_e[2] & input_d[1]);
  assign cgp_core_032 = ~(input_c[1] ^ input_a[1]);
  assign cgp_core_033_not = ~input_d[1];
  assign cgp_core_034 = ~input_c[1];
  assign cgp_core_035 = input_a[1] & input_b[1];
  assign cgp_core_036 = input_b[2] ^ cgp_core_026;
  assign cgp_core_037 = input_b[2] & cgp_core_026;
  assign cgp_core_038 = cgp_core_036 ^ cgp_core_035;
  assign cgp_core_039 = cgp_core_036 & cgp_core_035;
  assign cgp_core_040 = cgp_core_037 | cgp_core_039;
  assign cgp_core_044 = ~(input_d[2] | input_d[0]);
  assign cgp_core_045_not = ~input_e[0];
  assign cgp_core_050 = input_a[2] ^ input_d[2];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_052 = cgp_core_050 ^ input_a[1];
  assign cgp_core_053 = cgp_core_050 & input_a[1];
  assign cgp_core_054 = cgp_core_051 | cgp_core_053;
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_057 = cgp_core_040 & cgp_core_056;
  assign cgp_core_059 = ~(cgp_core_040 ^ cgp_core_054);
  assign cgp_core_061 = ~(input_c[0] | input_e[0]);
  assign cgp_core_063 = cgp_core_038 & cgp_core_059;
  assign cgp_core_064_not = ~cgp_core_052;
  assign cgp_core_065 = cgp_core_064_not & cgp_core_059;
  assign cgp_core_067 = ~(input_d[2] ^ input_a[1]);
  assign cgp_core_069 = input_e[0] | input_c[1];
  assign cgp_core_071 = input_c[2] ^ input_d[0];
  assign cgp_core_074_not = ~input_a[1];
  assign cgp_core_075 = input_a[1] ^ input_d[2];
  assign cgp_core_076 = cgp_core_065 | cgp_core_063;
  assign cgp_core_079 = cgp_core_057 | cgp_core_025;
  assign cgp_core_080 = cgp_core_076 | cgp_core_079;

  assign cgp_out[0] = cgp_core_080;
endmodule