module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_076;

  assign cgp_core_017 = input_b[1] & input_d[0];
  assign cgp_core_018 = input_c[0] ^ input_d[1];
  assign cgp_core_021 = ~(input_c[1] & input_b[0]);
  assign cgp_core_022 = ~input_a[2];
  assign cgp_core_024 = input_b[2] ^ input_e[1];
  assign cgp_core_025 = ~(input_b[2] ^ input_c[2]);
  assign cgp_core_026 = ~input_d[0];
  assign cgp_core_028_not = ~input_c[1];
  assign cgp_core_029 = input_b[2] ^ input_a[0];
  assign cgp_core_030 = ~(input_d[0] | input_e[1]);
  assign cgp_core_031 = input_b[2] | input_a[2];
  assign cgp_core_033 = input_d[0] | cgp_core_030;
  assign cgp_core_034 = ~(input_e[0] ^ input_a[2]);
  assign cgp_core_039 = ~input_e[1];
  assign cgp_core_041 = ~(input_c[0] ^ input_b[1]);
  assign cgp_core_043 = cgp_core_021 | input_a[1];
  assign cgp_core_044 = input_c[2] ^ input_a[2];
  assign cgp_core_047 = ~input_d[1];
  assign cgp_core_051 = input_b[2] ^ input_a[0];
  assign cgp_core_052 = ~(input_a[1] & input_d[2]);
  assign cgp_core_059 = ~input_d[2];
  assign cgp_core_060 = input_a[2] ^ input_e[2];
  assign cgp_core_061 = ~input_c[0];
  assign cgp_core_062 = input_d[2] | input_e[2];
  assign cgp_core_065 = ~input_e[1];
  assign cgp_core_069 = input_d[0] & input_a[1];
  assign cgp_core_070 = ~input_b[1];
  assign cgp_core_072 = input_b[1] | input_c[0];
  assign cgp_core_076 = ~(input_b[2] ^ input_b[1]);

  assign cgp_out[0] = 1'b0;
endmodule