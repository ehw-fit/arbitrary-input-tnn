module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059_not;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = input_g[0] & input_g[1];
  assign cgp_core_017 = ~(input_e[1] ^ input_f[0]);
  assign cgp_core_018 = ~(input_e[1] ^ input_g[1]);
  assign cgp_core_019 = input_e[1] & input_d[1];
  assign cgp_core_020 = input_e[0] | input_a[0];
  assign cgp_core_021_not = ~input_g[1];
  assign cgp_core_023 = ~(input_b[0] | input_a[1]);
  assign cgp_core_024 = input_a[1] | input_g[1];
  assign cgp_core_026 = input_a[1] & cgp_core_020;
  assign cgp_core_028 = input_e[1] & input_e[1];
  assign cgp_core_030 = ~input_g[1];
  assign cgp_core_031 = ~(cgp_core_019 | cgp_core_026);
  assign cgp_core_033 = ~(input_g[0] & input_a[1]);
  assign cgp_core_034 = ~(input_b[1] | input_b[1]);
  assign cgp_core_036 = input_b[1] ^ input_d[1];
  assign cgp_core_037_not = ~input_c[1];
  assign cgp_core_038 = input_c[0] | input_e[0];
  assign cgp_core_039 = input_e[0] ^ input_g[1];
  assign cgp_core_040 = ~(input_g[1] ^ input_d[1]);
  assign cgp_core_041 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_044 = ~(input_a[0] | input_b[0]);
  assign cgp_core_045 = input_c[1] ^ input_a[1];
  assign cgp_core_046 = ~input_c[1];
  assign cgp_core_047 = ~(input_e[0] & input_a[0]);
  assign cgp_core_048 = ~(input_a[1] & input_g[0]);
  assign cgp_core_050 = ~(input_c[0] & input_f[1]);
  assign cgp_core_051 = ~(input_a[1] | input_b[0]);
  assign cgp_core_052 = ~input_c[0];
  assign cgp_core_054 = input_b[1] & input_f[1];
  assign cgp_core_055 = ~(input_a[0] | input_e[1]);
  assign cgp_core_056 = input_c[1] & input_g[1];
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058 = input_d[0] & input_d[0];
  assign cgp_core_059_not = ~input_e[1];
  assign cgp_core_060 = ~(cgp_core_031 | cgp_core_057);
  assign cgp_core_063 = ~(input_e[1] ^ input_g[1]);
  assign cgp_core_066 = ~(input_d[0] | input_a[0]);
  assign cgp_core_067 = input_c[0] | input_g[0];
  assign cgp_core_068 = input_b[0] | input_a[0];
  assign cgp_core_070 = ~(input_f[0] | input_b[1]);
  assign cgp_core_071 = ~(input_f[1] | input_a[0]);
  assign cgp_core_075 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_076 = ~(input_f[0] & input_b[1]);
  assign cgp_core_077 = input_f[0] ^ input_f[0];
  assign cgp_core_078 = ~(input_c[1] | input_f[0]);
  assign cgp_core_079 = input_a[0] & input_g[0];

  assign cgp_out[0] = cgp_core_060;
endmodule