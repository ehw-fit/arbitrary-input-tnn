module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_067_not;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081_not;
  wire cgp_core_082;
  wire cgp_core_083;

  assign cgp_core_016 = ~(input_g[0] | input_g[1]);
  assign cgp_core_017 = input_c[0] & input_a[0];
  assign cgp_core_018 = input_a[1] | input_c[1];
  assign cgp_core_019 = input_a[1] & input_c[1];
  assign cgp_core_020 = cgp_core_018 | cgp_core_017;
  assign cgp_core_021 = cgp_core_018 & cgp_core_017;
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_024 = input_g[0] | input_e[0];
  assign cgp_core_026 = input_g[0] & input_a[0];
  assign cgp_core_028 = ~(input_d[0] & input_c[0]);
  assign cgp_core_029 = input_d[1] | input_c[0];
  assign cgp_core_030 = ~(input_d[1] | input_g[1]);
  assign cgp_core_032 = input_d[1] | input_e[1];
  assign cgp_core_033 = input_d[1] & input_e[1];
  assign cgp_core_035 = ~input_f[1];
  assign cgp_core_037 = input_g[1] | cgp_core_033;
  assign cgp_core_039 = ~(input_d[1] & input_g[0]);
  assign cgp_core_040_not = ~input_d[1];
  assign cgp_core_041 = cgp_core_020 | cgp_core_032;
  assign cgp_core_042 = cgp_core_020 & cgp_core_032;
  assign cgp_core_043 = cgp_core_041 | input_g[0];
  assign cgp_core_046 = cgp_core_022 | cgp_core_037;
  assign cgp_core_047 = input_b[0] & input_a[1];
  assign cgp_core_048 = cgp_core_046 | cgp_core_042;
  assign cgp_core_051 = ~(input_e[1] ^ input_g[1]);
  assign cgp_core_052 = ~(input_a[0] ^ input_e[1]);
  assign cgp_core_053_not = ~input_a[0];
  assign cgp_core_054 = input_c[1] & input_c[1];
  assign cgp_core_056 = input_b[1] & input_f[1];
  assign cgp_core_060 = input_d[0] ^ input_c[1];
  assign cgp_core_061 = input_a[1] & input_g[1];
  assign cgp_core_062 = input_d[1] & input_f[1];
  assign cgp_core_067_not = ~cgp_core_056;
  assign cgp_core_071 = cgp_core_043 & cgp_core_067_not;
  assign cgp_core_072 = ~(input_g[1] ^ input_b[1]);
  assign cgp_core_073 = input_f[0] & input_d[1];
  assign cgp_core_076 = ~(input_f[1] & input_d[0]);
  assign cgp_core_078 = input_e[0] ^ input_a[1];
  assign cgp_core_079 = cgp_core_071 | cgp_core_048;
  assign cgp_core_081_not = ~input_c[0];
  assign cgp_core_082 = ~(input_a[1] ^ input_g[0]);
  assign cgp_core_083 = input_c[1] | input_g[1];

  assign cgp_out[0] = cgp_core_079;
endmodule