module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068_not;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_080_not;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;

  assign cgp_core_021 = input_f[1] ^ input_f[1];
  assign cgp_core_022 = ~input_h[0];
  assign cgp_core_023 = input_f[1] & input_h[1];
  assign cgp_core_024 = input_e[1] | input_g[0];
  assign cgp_core_026 = input_a[1] & input_e[0];
  assign cgp_core_027 = input_e[0] | input_g[0];
  assign cgp_core_028 = input_a[1] & input_a[1];
  assign cgp_core_029 = ~(input_g[1] | input_b[0]);
  assign cgp_core_030 = ~input_b[1];
  assign cgp_core_031 = ~input_a[0];
  assign cgp_core_032 = input_h[0] ^ input_e[1];
  assign cgp_core_034 = ~(input_g[0] | input_b[1]);
  assign cgp_core_035 = input_c[0] & input_a[0];
  assign cgp_core_036 = input_f[1] & input_c[0];
  assign cgp_core_037 = input_g[1] & input_b[0];
  assign cgp_core_038 = ~(input_h[1] | input_b[0]);
  assign cgp_core_039 = ~(input_g[1] | input_f[1]);
  assign cgp_core_040 = input_g[1] | input_g[1];
  assign cgp_core_041 = input_d[1] & cgp_core_034;
  assign cgp_core_047 = ~(input_f[0] & input_e[0]);
  assign cgp_core_048 = input_e[1] ^ input_a[0];
  assign cgp_core_049 = input_g[0] | input_b[1];
  assign cgp_core_050 = ~(input_c[1] & input_c[1]);
  assign cgp_core_051 = input_a[0] & cgp_core_041;
  assign cgp_core_052 = cgp_core_029 ^ input_g[0];
  assign cgp_core_054_not = ~input_d[0];
  assign cgp_core_055 = ~cgp_core_052;
  assign cgp_core_061 = ~(input_c[0] ^ input_a[1]);
  assign cgp_core_062 = input_b[0] & input_b[0];
  assign cgp_core_065 = input_h[0] & input_f[0];
  assign cgp_core_067 = ~(input_e[0] | input_c[0]);
  assign cgp_core_068_not = ~input_h[1];
  assign cgp_core_069_not = ~input_f[0];
  assign cgp_core_070 = ~input_e[0];
  assign cgp_core_071 = ~(input_f[1] | input_h[0]);
  assign cgp_core_072 = input_a[1] & input_f[1];
  assign cgp_core_073 = cgp_core_070 & input_h[0];
  assign cgp_core_080_not = ~input_h[1];
  assign cgp_core_081 = ~(input_b[1] ^ input_g[0]);
  assign cgp_core_082 = input_c[0] ^ input_d[0];
  assign cgp_core_084 = input_c[1] & input_a[0];
  assign cgp_core_085 = ~(cgp_core_084 ^ cgp_core_082);
  assign cgp_core_086 = ~(cgp_core_054_not | input_a[1]);
  assign cgp_core_088 = input_e[0] ^ input_b[1];
  assign cgp_core_089 = cgp_core_050 & cgp_core_088;
  assign cgp_core_091 = ~(input_b[0] ^ input_g[1]);
  assign cgp_core_092 = input_f[0] ^ input_a[1];
  assign cgp_core_093 = input_e[1] | input_f[1];
  assign cgp_core_094 = input_h[0] | input_c[1];

  assign cgp_out[0] = 1'b1;
endmodule