module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_082;
  wire cgp_core_083;

  assign cgp_core_016_not = ~input_g[1];
  assign cgp_core_017 = ~(input_g[1] ^ input_f[1]);
  assign cgp_core_018 = ~(input_e[0] ^ input_f[1]);
  assign cgp_core_019 = ~(input_a[1] | input_b[0]);
  assign cgp_core_021 = ~(input_a[0] & input_b[0]);
  assign cgp_core_022 = input_f[1] | input_a[0];
  assign cgp_core_023 = ~(input_f[1] | input_b[0]);
  assign cgp_core_025 = ~input_e[0];
  assign cgp_core_026 = input_a[0] ^ input_d[0];
  assign cgp_core_027 = ~(input_g[1] & input_g[1]);
  assign cgp_core_028_not = ~input_f[0];
  assign cgp_core_029 = input_e[1] | input_a[1];
  assign cgp_core_032 = ~(input_c[1] | input_e[1]);
  assign cgp_core_033 = ~input_b[1];
  assign cgp_core_035 = input_a[1] & input_c[1];
  assign cgp_core_036 = input_d[0] | input_g[1];
  assign cgp_core_037 = cgp_core_029 | input_d[1];
  assign cgp_core_039 = ~(input_g[0] | input_b[0]);
  assign cgp_core_041 = ~input_c[1];
  assign cgp_core_043 = input_b[1] & input_c[1];
  assign cgp_core_044 = ~(input_c[1] & input_b[0]);
  assign cgp_core_046 = input_g[1] ^ input_a[1];
  assign cgp_core_048 = input_f[1] | input_b[1];
  assign cgp_core_051 = input_c[1] | cgp_core_037;
  assign cgp_core_053 = ~input_g[0];
  assign cgp_core_054_not = ~input_d[0];
  assign cgp_core_055 = ~input_f[1];
  assign cgp_core_056 = ~(input_f[1] & input_f[1]);
  assign cgp_core_057 = input_e[0] | input_b[0];
  assign cgp_core_060 = ~(input_g[1] & input_b[1]);
  assign cgp_core_062 = ~(input_c[0] ^ input_f[0]);
  assign cgp_core_063 = input_e[0] ^ input_d[1];
  assign cgp_core_066 = ~(input_f[1] | input_c[0]);
  assign cgp_core_069 = input_a[1] ^ input_e[0];
  assign cgp_core_071 = input_g[0] | input_d[1];
  assign cgp_core_072 = ~input_b[1];
  assign cgp_core_076 = input_f[1] | input_d[0];
  assign cgp_core_077 = input_a[0] & input_b[1];
  assign cgp_core_082 = cgp_core_051 | input_g[1];
  assign cgp_core_083 = ~(input_b[0] & input_b[0]);

  assign cgp_out[0] = cgp_core_082;
endmodule