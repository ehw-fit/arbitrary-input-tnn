module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055_not;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_079;
  wire cgp_core_080_not;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_094_not;

  assign cgp_core_018 = input_d[0] | input_c[1];
  assign cgp_core_019 = input_b[0] & input_a[1];
  assign cgp_core_021 = input_h[1] & input_c[1];
  assign cgp_core_027 = ~(input_c[0] | input_c[1]);
  assign cgp_core_028 = ~(input_h[0] & input_f[0]);
  assign cgp_core_029 = input_c[0] ^ input_g[1];
  assign cgp_core_030 = input_a[1] ^ input_a[0];
  assign cgp_core_031 = input_f[1] | input_b[1];
  assign cgp_core_033 = ~input_a[1];
  assign cgp_core_035 = ~(input_c[0] | input_h[1]);
  assign cgp_core_036 = input_g[1] & input_e[0];
  assign cgp_core_037 = input_d[1] ^ input_h[0];
  assign cgp_core_038 = ~(input_g[1] | input_f[1]);
  assign cgp_core_040 = input_a[1] ^ input_f[1];
  assign cgp_core_041 = ~input_h[1];
  assign cgp_core_042 = input_h[1] & input_h[0];
  assign cgp_core_043 = ~(input_d[1] ^ input_f[0]);
  assign cgp_core_044 = ~(input_g[0] & input_c[0]);
  assign cgp_core_045 = input_e[0] & input_f[0];
  assign cgp_core_046 = ~input_h[0];
  assign cgp_core_047 = ~(cgp_core_044 | input_h[0]);
  assign cgp_core_048 = ~input_a[1];
  assign cgp_core_049 = ~input_d[0];
  assign cgp_core_050 = input_a[0] & input_d[1];
  assign cgp_core_052 = cgp_core_029 & cgp_core_045;
  assign cgp_core_054 = ~input_b[0];
  assign cgp_core_055_not = ~cgp_core_052;
  assign cgp_core_056 = ~(input_b[1] | input_d[0]);
  assign cgp_core_059 = input_f[1] & input_g[1];
  assign cgp_core_061 = ~(input_e[0] & input_a[0]);
  assign cgp_core_062 = ~input_a[0];
  assign cgp_core_064 = input_e[1] | input_a[0];
  assign cgp_core_067 = input_h[1] & input_f[0];
  assign cgp_core_068 = ~(input_a[0] | input_e[0]);
  assign cgp_core_070 = ~(input_b[1] | input_c[0]);
  assign cgp_core_071 = ~(input_b[1] | input_e[0]);
  assign cgp_core_072 = ~(input_g[0] ^ input_b[1]);
  assign cgp_core_073 = input_e[0] | input_b[1];
  assign cgp_core_074 = input_c[0] ^ input_e[0];
  assign cgp_core_076 = input_b[0] | cgp_core_064;
  assign cgp_core_079 = ~(input_f[0] ^ input_d[1]);
  assign cgp_core_080_not = ~input_e[1];
  assign cgp_core_081 = cgp_core_059 | input_a[0];
  assign cgp_core_082 = ~input_f[0];
  assign cgp_core_083 = ~(input_g[0] ^ input_e[0]);
  assign cgp_core_084 = input_b[0] & input_e[0];
  assign cgp_core_085 = ~input_c[0];
  assign cgp_core_086 = ~input_b[0];
  assign cgp_core_088 = ~(input_d[1] ^ input_b[1]);
  assign cgp_core_089 = ~(input_f[0] ^ input_e[0]);
  assign cgp_core_094_not = ~input_h[0];

  assign cgp_out[0] = 1'b1;
endmodule