module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_039_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075_not;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;

  assign cgp_core_019 = ~(input_a[13] & input_a[7]);
  assign cgp_core_021 = input_a[11] ^ input_a[10];
  assign cgp_core_022 = input_a[8] | input_a[13];
  assign cgp_core_023 = input_a[2] | input_a[5];
  assign cgp_core_024 = ~(input_a[7] ^ input_a[3]);
  assign cgp_core_025_not = ~input_a[11];
  assign cgp_core_027 = ~(input_a[5] | input_a[1]);
  assign cgp_core_030 = input_a[0] ^ input_a[4];
  assign cgp_core_032 = input_a[13] & input_a[3];
  assign cgp_core_033 = input_a[13] | input_a[5];
  assign cgp_core_035_not = ~input_a[13];
  assign cgp_core_036 = ~input_a[2];
  assign cgp_core_037_not = ~input_a[7];
  assign cgp_core_039_not = ~input_a[12];
  assign cgp_core_041 = input_a[4] & input_a[8];
  assign cgp_core_042 = ~input_a[1];
  assign cgp_core_043 = input_a[2] ^ input_a[7];
  assign cgp_core_044 = ~input_a[4];
  assign cgp_core_046 = ~input_a[12];
  assign cgp_core_047 = input_a[0] ^ input_a[0];
  assign cgp_core_051 = ~(input_a[4] | input_a[0]);
  assign cgp_core_052 = input_a[0] ^ input_a[6];
  assign cgp_core_055 = ~input_a[5];
  assign cgp_core_058 = ~(input_a[4] ^ input_a[1]);
  assign cgp_core_060 = ~input_a[10];
  assign cgp_core_061 = ~(input_a[9] & input_a[7]);
  assign cgp_core_064 = ~(input_a[8] ^ input_a[12]);
  assign cgp_core_067 = ~(input_a[12] ^ input_a[3]);
  assign cgp_core_070 = ~input_a[7];
  assign cgp_core_071 = input_a[12] ^ input_a[9];
  assign cgp_core_072 = ~(input_a[9] ^ input_a[4]);
  assign cgp_core_073 = input_a[11] | input_a[0];
  assign cgp_core_074 = ~(input_a[4] ^ input_a[4]);
  assign cgp_core_075_not = ~input_a[12];
  assign cgp_core_076 = ~(input_a[12] ^ input_a[13]);
  assign cgp_core_077 = ~input_a[0];
  assign cgp_core_080 = input_a[7] & input_a[9];
  assign cgp_core_081 = ~(input_a[9] & input_a[6]);
  assign cgp_core_082 = input_a[7] ^ input_a[0];
  assign cgp_core_083 = ~(input_a[5] & input_a[12]);
  assign cgp_core_084 = ~(input_a[10] ^ input_a[7]);
  assign cgp_core_085 = ~(input_a[10] | input_a[4]);
  assign cgp_core_087 = input_a[1] ^ input_a[8];
  assign cgp_core_089 = ~input_a[5];
  assign cgp_core_090 = ~input_a[8];

  assign cgp_out[0] = input_a[9];
  assign cgp_out[1] = cgp_core_061;
  assign cgp_out[2] = cgp_core_061;
  assign cgp_out[3] = cgp_core_080;
endmodule