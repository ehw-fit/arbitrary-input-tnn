module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017 = ~(input_d[1] & input_c[0]);
  assign cgp_core_018 = input_d[2] ^ input_d[2];
  assign cgp_core_019 = input_b[0] ^ input_c[2];
  assign cgp_core_020 = ~input_c[0];
  assign cgp_core_023 = input_d[2] | input_b[1];
  assign cgp_core_025 = input_a[2] & input_b[2];
  assign cgp_core_026 = ~(input_e[0] & input_d[2]);
  assign cgp_core_027 = input_a[2] & input_a[1];
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_032 = ~input_c[0];
  assign cgp_core_034 = ~(input_d[2] & input_e[0]);
  assign cgp_core_036 = input_a[2] | input_e[0];
  assign cgp_core_039 = input_d[2] & input_c[2];
  assign cgp_core_044 = ~(input_a[0] ^ input_b[2]);
  assign cgp_core_047 = input_d[2] | input_c[2];
  assign cgp_core_048 = ~(input_a[1] | input_d[1]);
  assign cgp_core_049 = ~(input_c[1] ^ input_c[0]);
  assign cgp_core_050 = ~input_e[0];
  assign cgp_core_051 = input_e[2] & cgp_core_047;
  assign cgp_core_053 = cgp_core_039 | cgp_core_051;
  assign cgp_core_054 = input_a[0] ^ input_c[0];
  assign cgp_core_055 = ~(input_d[1] & input_e[1]);
  assign cgp_core_057 = ~cgp_core_053;
  assign cgp_core_058 = cgp_core_028 & cgp_core_057;
  assign cgp_core_059 = input_e[0] ^ input_c[0];
  assign cgp_core_062 = input_c[0] ^ input_b[1];
  assign cgp_core_063 = ~(input_b[0] ^ input_d[2]);
  assign cgp_core_064 = input_a[2] & input_a[0];
  assign cgp_core_066 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_068 = input_a[0] | input_b[2];
  assign cgp_core_070 = ~(input_d[0] ^ input_c[2]);
  assign cgp_core_073 = input_a[2] ^ input_d[1];
  assign cgp_core_074 = ~(input_e[0] ^ input_e[0]);
  assign cgp_core_076 = ~(input_b[2] | input_c[0]);
  assign cgp_core_077 = ~(input_d[1] & input_c[1]);
  assign cgp_core_079 = ~(input_c[2] & input_b[0]);
  assign cgp_core_080 = ~(input_e[0] & input_e[2]);

  assign cgp_out[0] = cgp_core_058;
endmodule