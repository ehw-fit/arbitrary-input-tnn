module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_043;
  wire cgp_core_046_not;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068_not;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_077;
  wire cgp_core_080;
  wire cgp_core_082_not;
  wire cgp_core_083;

  assign cgp_core_016 = input_a[0] ^ input_b[0];
  assign cgp_core_023 = ~(input_e[0] & input_g[0]);
  assign cgp_core_025 = input_e[1] ^ input_g[1];
  assign cgp_core_027 = cgp_core_025 | input_e[0];
  assign cgp_core_028 = cgp_core_025 | input_e[0];
  assign cgp_core_029 = input_a[1] | cgp_core_028;
  assign cgp_core_032 = input_d[1] ^ cgp_core_027;
  assign cgp_core_033 = input_d[0] ^ input_d[0];
  assign cgp_core_034_not = ~cgp_core_032;
  assign cgp_core_038 = cgp_core_029 & input_f[0];
  assign cgp_core_039 = cgp_core_016 ^ input_f[1];
  assign cgp_core_043 = ~input_d[1];
  assign cgp_core_046_not = ~input_d[0];
  assign cgp_core_050 = input_e[1] | input_b[1];
  assign cgp_core_053 = input_b[0] ^ input_g[0];
  assign cgp_core_054 = input_b[0] & input_f[0];
  assign cgp_core_055 = ~(input_b[1] ^ input_f[1]);
  assign cgp_core_057 = cgp_core_055 ^ input_d[1];
  assign cgp_core_058 = ~input_e[1];
  assign cgp_core_059 = ~(input_b[1] | cgp_core_058);
  assign cgp_core_064 = cgp_core_059 ^ input_e[1];
  assign cgp_core_067 = ~(input_a[0] & input_e[0]);
  assign cgp_core_068_not = ~input_f[1];
  assign cgp_core_069 = cgp_core_057 | cgp_core_057;
  assign cgp_core_070 = ~(cgp_core_043 | input_e[0]);
  assign cgp_core_071 = input_g[1] & cgp_core_068_not;
  assign cgp_core_072 = ~(cgp_core_043 ^ input_e[1]);
  assign cgp_core_074 = ~cgp_core_053;
  assign cgp_core_077 = ~(input_c[1] ^ input_c[1]);
  assign cgp_core_080 = input_b[0] | input_g[1];
  assign cgp_core_082_not = ~input_e[0];
  assign cgp_core_083 = input_a[1] | input_f[0];

  assign cgp_out[0] = 1'b1;
endmodule