module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_046_not;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_059;

  assign cgp_core_015 = ~(input_b[0] ^ input_d[2]);
  assign cgp_core_018 = ~(input_a[2] | input_a[0]);
  assign cgp_core_019 = ~(input_a[1] ^ input_a[2]);
  assign cgp_core_020 = ~(input_a[1] | input_c[0]);
  assign cgp_core_022_not = ~input_c[0];
  assign cgp_core_023 = input_d[2] | input_d[0];
  assign cgp_core_024 = input_c[1] & input_d[1];
  assign cgp_core_025 = ~(input_a[1] | input_a[1]);
  assign cgp_core_027 = ~(input_a[1] ^ input_c[2]);
  assign cgp_core_029 = ~(input_b[2] & input_b[0]);
  assign cgp_core_030 = ~(input_d[2] ^ input_c[2]);
  assign cgp_core_032 = ~(input_b[1] & input_b[2]);
  assign cgp_core_037 = input_a[1] & input_b[1];
  assign cgp_core_038 = ~(input_c[2] | input_c[1]);
  assign cgp_core_041 = ~input_c[2];
  assign cgp_core_042 = input_b[2] & cgp_core_041;
  assign cgp_core_046_not = ~input_c[2];
  assign cgp_core_048 = ~(input_a[0] | input_d[2]);
  assign cgp_core_049 = ~(input_a[1] | input_c[1]);
  assign cgp_core_052 = ~(input_d[2] | input_d[2]);
  assign cgp_core_053 = input_b[1] & input_c[0];
  assign cgp_core_054 = ~(input_b[0] & input_b[0]);
  assign cgp_core_056 = ~input_c[2];
  assign cgp_core_059 = input_a[2] | cgp_core_042;

  assign cgp_out[0] = cgp_core_059;
endmodule