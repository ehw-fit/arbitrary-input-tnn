module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_021 = ~input_b[2];
  assign cgp_core_023 = ~input_a[0];
  assign cgp_core_024 = input_e[2] | input_c[1];
  assign cgp_core_026 = ~(input_d[0] ^ input_a[2]);
  assign cgp_core_027 = input_c[1] & input_b[2];
  assign cgp_core_028 = input_c[2] & input_e[2];
  assign cgp_core_029 = input_c[0] & input_b[2];
  assign cgp_core_030 = input_d[1] | input_f[2];
  assign cgp_core_032 = input_d[0] & input_d[1];
  assign cgp_core_033 = input_d[1] & input_e[0];
  assign cgp_core_036 = input_e[2] ^ input_b[1];
  assign cgp_core_038 = input_e[0] ^ input_b[0];
  assign cgp_core_039 = ~(input_a[2] ^ input_e[2]);
  assign cgp_core_040 = ~(input_c[2] | input_e[2]);
  assign cgp_core_042 = ~input_d[2];
  assign cgp_core_043 = input_a[2] | input_c[2];
  assign cgp_core_044 = input_e[2] | cgp_core_043;
  assign cgp_core_045 = cgp_core_028 & input_a[2];
  assign cgp_core_046 = input_e[0] ^ input_e[0];
  assign cgp_core_047 = input_e[0] ^ input_a[0];
  assign cgp_core_048 = input_a[0] | input_b[0];
  assign cgp_core_049 = ~(input_b[2] | input_f[0]);
  assign cgp_core_050 = input_f[0] | input_f[0];
  assign cgp_core_051 = ~input_b[2];
  assign cgp_core_053 = input_d[2] | input_f[2];
  assign cgp_core_054 = input_d[2] & input_f[2];
  assign cgp_core_058 = ~input_d[2];
  assign cgp_core_059 = ~(input_f[1] | input_c[2]);
  assign cgp_core_061 = input_d[0] ^ input_b[1];
  assign cgp_core_062 = ~(input_a[2] & input_b[1]);
  assign cgp_core_063 = ~(input_d[2] & input_e[2]);
  assign cgp_core_064 = ~(input_a[0] ^ input_b[0]);
  assign cgp_core_065 = input_c[2] & input_d[1];
  assign cgp_core_066 = input_b[2] & cgp_core_053;
  assign cgp_core_068 = input_d[0] & input_b[2];
  assign cgp_core_070 = cgp_core_054 | cgp_core_066;
  assign cgp_core_071 = ~(input_f[1] & input_b[2]);
  assign cgp_core_072 = input_e[0] | input_c[2];
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = cgp_core_044 & cgp_core_075;
  assign cgp_core_078 = input_a[0] | input_d[2];
  assign cgp_core_079 = ~input_e[0];
  assign cgp_core_081 = ~(input_f[1] & input_e[0]);
  assign cgp_core_082 = input_f[2] | input_c[0];
  assign cgp_core_083 = input_e[1] | input_b[1];
  assign cgp_core_084 = ~input_f[2];
  assign cgp_core_085 = input_d[2] & input_a[1];
  assign cgp_core_086 = input_b[2] ^ input_f[2];
  assign cgp_core_088 = input_a[0] | input_e[2];
  assign cgp_core_089 = ~input_d[0];
  assign cgp_core_098 = cgp_core_076 | cgp_core_045;
  assign cgp_core_099 = input_b[1] & input_f[2];

  assign cgp_out[0] = cgp_core_098;
endmodule