module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_016 = input_c[0] ^ input_g[0];
  assign cgp_core_018 = input_f[1] | input_c[0];
  assign cgp_core_019 = ~input_b[1];
  assign cgp_core_022 = input_c[1] & input_d[0];
  assign cgp_core_026_not = ~input_d[0];
  assign cgp_core_027 = input_a[1] & input_b[1];
  assign cgp_core_029 = ~(input_b[1] | input_c[0]);
  assign cgp_core_030 = input_a[0] & input_e[1];
  assign cgp_core_031 = ~input_c[0];
  assign cgp_core_032 = input_f[1] & input_g[0];
  assign cgp_core_034 = ~(input_e[1] ^ input_d[0]);
  assign cgp_core_038 = input_c[0] & input_e[0];
  assign cgp_core_040 = input_c[0] & input_g[0];
  assign cgp_core_041 = input_g[1] | cgp_core_040;
  assign cgp_core_042 = ~(input_g[1] | input_c[0]);
  assign cgp_core_043 = ~(input_a[1] | input_b[1]);
  assign cgp_core_044 = input_b[0] | input_d[1];
  assign cgp_core_045 = ~input_e[1];
  assign cgp_core_047 = ~(input_e[0] & input_b[1]);
  assign cgp_core_049 = ~(input_f[0] ^ input_f[0]);
  assign cgp_core_050 = input_d[0] | input_b[1];
  assign cgp_core_052 = input_c[1] ^ input_g[1];
  assign cgp_core_053 = input_b[0] ^ input_c[1];
  assign cgp_core_054 = ~(input_f[1] & input_b[0]);
  assign cgp_core_055 = ~(input_g[1] ^ input_c[0]);
  assign cgp_core_057 = input_a[1] & input_f[1];
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = cgp_core_041 & cgp_core_058;
  assign cgp_core_061 = ~input_b[1];
  assign cgp_core_062 = input_d[1] & cgp_core_061;
  assign cgp_core_065 = input_b[1] & input_e[1];
  assign cgp_core_066 = input_b[1] | input_e[0];
  assign cgp_core_067 = ~(input_e[1] | input_c[0]);
  assign cgp_core_068 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_069 = ~(input_g[1] ^ input_a[0]);
  assign cgp_core_070 = input_e[0] & input_e[1];
  assign cgp_core_072 = input_c[0] | input_d[1];
  assign cgp_core_075 = input_c[1] & input_e[1];
  assign cgp_core_077 = cgp_core_059 | cgp_core_075;
  assign cgp_core_078 = cgp_core_062 | cgp_core_077;

  assign cgp_out[0] = cgp_core_078;
endmodule