module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_026_not;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_034_not;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_058_not;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_018 = input_c[1] ^ input_e[1];
  assign cgp_core_026_not = ~input_a[1];
  assign cgp_core_029 = input_b[0] | input_g[1];
  assign cgp_core_032 = ~(input_d[0] | input_a[0]);
  assign cgp_core_034_not = ~input_d[1];
  assign cgp_core_036 = input_b[1] ^ input_e[0];
  assign cgp_core_039 = input_g[0] ^ input_g[0];
  assign cgp_core_040 = input_d[1] & input_b[1];
  assign cgp_core_042 = ~(input_f[1] & input_g[1]);
  assign cgp_core_043 = ~(input_e[1] ^ input_a[0]);
  assign cgp_core_045 = input_c[0] | input_e[0];
  assign cgp_core_046 = input_c[0] ^ cgp_core_039;
  assign cgp_core_047 = input_e[0] & input_g[1];
  assign cgp_core_048 = ~(input_a[0] & cgp_core_043);
  assign cgp_core_049 = cgp_core_036 ^ input_c[0];
  assign cgp_core_050 = ~(cgp_core_048 | input_d[1]);
  assign cgp_core_052 = ~input_a[1];
  assign cgp_core_058_not = ~input_g[0];
  assign cgp_core_059 = input_e[0] & cgp_core_058_not;
  assign cgp_core_060 = ~(input_a[0] ^ input_d[1]);
  assign cgp_core_061 = ~input_a[1];
  assign cgp_core_066 = ~(cgp_core_050 & input_f[0]);
  assign cgp_core_067 = input_g[0] & cgp_core_066;
  assign cgp_core_068 = input_a[0] & input_f[1];
  assign cgp_core_069 = ~(input_f[0] ^ input_f[0]);
  assign cgp_core_071 = ~input_e[0];
  assign cgp_core_072 = input_f[0] ^ input_b[0];
  assign cgp_core_073 = ~(cgp_core_072 & input_f[1]);
  assign cgp_core_074 = ~(input_c[0] ^ cgp_core_046);
  assign cgp_core_076 = ~(input_g[1] ^ input_g[0]);
  assign cgp_core_077 = input_b[1] | input_f[0];
  assign cgp_core_078 = input_b[0] | input_b[0];
  assign cgp_core_079 = cgp_core_076 | input_b[0];

  assign cgp_out[0] = input_e[0];
endmodule