module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056_not;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_080;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_097;

  assign cgp_core_020 = input_d[2] ^ input_c[1];
  assign cgp_core_021 = ~(input_b[2] ^ input_f[1]);
  assign cgp_core_022 = ~(input_a[1] | input_c[0]);
  assign cgp_core_024 = input_f[2] ^ input_b[1];
  assign cgp_core_027 = input_a[2] ^ input_b[2];
  assign cgp_core_028 = input_a[2] ^ input_b[2];
  assign cgp_core_034 = ~(input_b[1] | input_f[2]);
  assign cgp_core_037 = ~(input_c[2] ^ input_b[1]);
  assign cgp_core_041 = input_f[2] ^ input_a[2];
  assign cgp_core_044 = ~input_d[2];
  assign cgp_core_045 = input_a[1] | input_a[0];
  assign cgp_core_046 = ~(input_e[0] ^ input_f[1]);
  assign cgp_core_047 = input_c[1] & input_f[1];
  assign cgp_core_048 = input_b[0] ^ input_f[0];
  assign cgp_core_049 = cgp_core_046 | cgp_core_045;
  assign cgp_core_050 = ~input_c[2];
  assign cgp_core_052 = input_b[2] & input_f[0];
  assign cgp_core_053 = ~(input_a[0] & cgp_core_050);
  assign cgp_core_054 = ~(input_a[2] ^ input_c[0]);
  assign cgp_core_055 = cgp_core_052 ^ input_d[0];
  assign cgp_core_056_not = ~input_e[2];
  assign cgp_core_057 = input_d[0] & cgp_core_044;
  assign cgp_core_058 = input_a[1] & cgp_core_048;
  assign cgp_core_061 = input_b[1] & input_e[1];
  assign cgp_core_062 = input_b[2] | cgp_core_061;
  assign cgp_core_064 = cgp_core_041 ^ cgp_core_053;
  assign cgp_core_065 = input_b[0] | input_d[0];
  assign cgp_core_066 = ~(input_f[1] & input_b[1]);
  assign cgp_core_067 = cgp_core_064 & input_a[2];
  assign cgp_core_068 = ~(input_a[2] & cgp_core_055);
  assign cgp_core_070 = ~(input_f[1] ^ input_b[1]);
  assign cgp_core_071 = ~input_a[2];
  assign cgp_core_072 = ~(cgp_core_055 & input_b[1]);
  assign cgp_core_073 = ~(cgp_core_072 & input_b[1]);
  assign cgp_core_074 = input_f[1] | input_d[2];
  assign cgp_core_076 = input_f[1] & input_c[1];
  assign cgp_core_077 = input_f[0] & input_d[1];
  assign cgp_core_080 = ~input_d[0];
  assign cgp_core_084 = ~(input_f[0] | input_e[1]);
  assign cgp_core_085 = ~input_b[2];
  assign cgp_core_086 = ~(cgp_core_024 | input_f[1]);
  assign cgp_core_087 = ~(input_e[2] ^ input_e[2]);
  assign cgp_core_089 = ~input_a[1];
  assign cgp_core_092 = ~(input_e[2] ^ input_b[1]);
  assign cgp_core_093 = ~(input_b[1] | input_d[1]);
  assign cgp_core_094 = ~cgp_core_093;
  assign cgp_core_095 = cgp_core_087 | input_b[1];
  assign cgp_core_097 = cgp_core_077 | cgp_core_094;

  assign cgp_out[0] = 1'b0;
endmodule