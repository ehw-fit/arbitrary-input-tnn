module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;

  assign cgp_core_021 = input_f[1] & input_e[1];
  assign cgp_core_022 = ~(input_b[0] ^ input_h[1]);
  assign cgp_core_025 = ~input_g[0];
  assign cgp_core_026 = ~input_g[1];
  assign cgp_core_028 = input_c[1] | input_f[1];
  assign cgp_core_030 = ~(input_h[1] | input_d[0]);
  assign cgp_core_032 = ~(input_f[0] & input_c[0]);
  assign cgp_core_033 = input_c[1] & input_g[1];
  assign cgp_core_035 = ~input_h[1];
  assign cgp_core_036 = ~(input_f[0] & input_c[1]);
  assign cgp_core_038 = ~(input_d[1] | input_c[1]);
  assign cgp_core_039 = input_d[0] & input_a[1];
  assign cgp_core_040 = input_a[0] | input_c[1];
  assign cgp_core_042 = ~(input_d[0] & input_g[0]);
  assign cgp_core_045 = ~input_d[0];
  assign cgp_core_047 = input_g[0] | input_b[1];
  assign cgp_core_049 = ~(input_h[1] & input_e[0]);
  assign cgp_core_050 = input_e[1] ^ input_a[0];
  assign cgp_core_051 = input_f[0] & input_g[0];
  assign cgp_core_052 = input_c[1] ^ input_f[0];
  assign cgp_core_054 = ~(input_h[0] | cgp_core_051);
  assign cgp_core_056 = ~(input_d[1] | input_a[1]);
  assign cgp_core_058 = ~input_g[1];
  assign cgp_core_059 = ~(input_f[1] | input_g[0]);
  assign cgp_core_062 = input_b[0] | input_e[0];
  assign cgp_core_063 = input_h[0] & cgp_core_049;
  assign cgp_core_067 = ~(input_d[0] & input_c[0]);
  assign cgp_core_068 = input_e[1] ^ input_c[1];
  assign cgp_core_076 = input_a[0] & input_h[0];
  assign cgp_core_078 = input_f[0] | input_c[0];
  assign cgp_core_080 = ~input_a[0];
  assign cgp_core_081 = input_h[0] ^ input_a[0];
  assign cgp_core_086 = ~(input_h[0] | input_f[1]);
  assign cgp_core_087 = ~(input_a[1] & input_h[1]);
  assign cgp_core_089 = input_f[0] & input_d[0];
  assign cgp_core_092 = ~input_g[0];
  assign cgp_core_093 = input_e[1] & input_a[1];
  assign cgp_core_094 = ~(input_d[1] & input_c[1]);
  assign cgp_core_095 = input_g[0] | input_d[0];

  assign cgp_out[0] = 1'b1;
endmodule