module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076_not;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_082;
  wire cgp_core_083;

  assign cgp_core_016 = input_e[1] | input_f[1];
  assign cgp_core_018 = input_a[1] | input_c[1];
  assign cgp_core_019 = input_a[1] & input_c[1];
  assign cgp_core_021 = input_a[0] | input_d[0];
  assign cgp_core_023 = ~input_e[1];
  assign cgp_core_024 = input_f[0] ^ input_g[1];
  assign cgp_core_025 = input_e[1] ^ input_g[1];
  assign cgp_core_026 = input_f[0] | input_g[1];
  assign cgp_core_027 = ~cgp_core_025;
  assign cgp_core_028 = ~(input_c[1] & input_g[1]);
  assign cgp_core_029 = input_g[1] | input_e[1];
  assign cgp_core_030 = ~(input_b[1] | input_d[0]);
  assign cgp_core_032 = input_d[1] ^ cgp_core_027;
  assign cgp_core_034 = cgp_core_032 ^ input_c[0];
  assign cgp_core_036 = input_d[1] | cgp_core_032;
  assign cgp_core_037 = cgp_core_029 | input_d[1];
  assign cgp_core_038 = cgp_core_029 & cgp_core_036;
  assign cgp_core_039 = input_a[0] | input_b[1];
  assign cgp_core_040 = ~(input_c[0] ^ input_g[1]);
  assign cgp_core_041 = cgp_core_018 ^ cgp_core_034;
  assign cgp_core_042 = cgp_core_018 & cgp_core_034;
  assign cgp_core_044 = input_g[0] & input_d[0];
  assign cgp_core_046 = input_c[0] | cgp_core_037;
  assign cgp_core_048 = cgp_core_046 | cgp_core_042;
  assign cgp_core_049 = input_c[0] & cgp_core_042;
  assign cgp_core_050 = cgp_core_019 | cgp_core_049;
  assign cgp_core_054 = input_f[0] & input_c[0];
  assign cgp_core_055 = input_b[1] ^ input_f[1];
  assign cgp_core_056 = input_b[1] & input_f[1];
  assign cgp_core_057 = cgp_core_055 ^ cgp_core_054;
  assign cgp_core_058 = cgp_core_055 & cgp_core_054;
  assign cgp_core_059 = cgp_core_056 | cgp_core_058;
  assign cgp_core_062 = ~input_d[1];
  assign cgp_core_064 = ~cgp_core_059;
  assign cgp_core_065 = cgp_core_048 & cgp_core_064;
  assign cgp_core_067 = ~(cgp_core_048 ^ cgp_core_059);
  assign cgp_core_069 = ~cgp_core_057;
  assign cgp_core_070 = cgp_core_041 & cgp_core_069;
  assign cgp_core_071 = cgp_core_070 & cgp_core_067;
  assign cgp_core_072 = ~(input_b[0] ^ input_e[1]);
  assign cgp_core_073 = input_b[0] ^ input_a[1];
  assign cgp_core_075 = input_b[0] | input_c[0];
  assign cgp_core_076_not = ~input_a[1];
  assign cgp_core_078 = input_a[1] | input_c[0];
  assign cgp_core_079 = cgp_core_071 | cgp_core_065;
  assign cgp_core_082 = cgp_core_050 | cgp_core_038;
  assign cgp_core_083 = cgp_core_079 | cgp_core_082;

  assign cgp_out[0] = cgp_core_083;
endmodule