module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_017 = input_a[1] & input_b[2];
  assign cgp_core_019 = input_e[0] ^ input_c[2];
  assign cgp_core_020 = ~(input_b[0] & input_d[0]);
  assign cgp_core_026 = ~(input_e[0] & input_c[2]);
  assign cgp_core_027 = input_e[2] & input_b[2];
  assign cgp_core_028_not = ~input_d[1];
  assign cgp_core_037 = input_a[1] ^ input_e[1];
  assign cgp_core_038 = ~(input_a[1] ^ input_b[0]);
  assign cgp_core_039 = ~(input_c[1] ^ input_b[0]);
  assign cgp_core_040 = input_a[2] & input_a[1];
  assign cgp_core_041 = input_a[2] ^ input_d[1];
  assign cgp_core_042 = ~(input_a[1] & input_a[2]);
  assign cgp_core_045 = ~input_c[0];
  assign cgp_core_046 = input_a[1] & input_c[0];
  assign cgp_core_049 = ~(input_c[2] | input_a[0]);
  assign cgp_core_050 = ~input_b[2];
  assign cgp_core_051 = input_c[1] | input_c[0];
  assign cgp_core_052 = ~input_c[0];
  assign cgp_core_054_not = ~input_d[0];
  assign cgp_core_055 = input_a[0] ^ input_d[2];
  assign cgp_core_058 = ~input_d[2];
  assign cgp_core_060 = input_d[2] ^ input_b[1];
  assign cgp_core_065 = ~input_c[0];
  assign cgp_core_066 = ~(input_d[0] & input_e[0]);
  assign cgp_core_068 = input_d[1] | input_a[2];
  assign cgp_core_069 = input_b[1] & input_c[2];
  assign cgp_core_071 = ~input_b[2];
  assign cgp_core_076 = ~input_b[0];
  assign cgp_core_077 = ~(input_e[1] & input_b[0]);
  assign cgp_core_079 = input_d[2] | input_b[2];

  assign cgp_out[0] = 1'b0;
endmodule