module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_058;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;

  assign cgp_core_014 = input_a[0] ^ input_c[0];
  assign cgp_core_015 = input_a[0] & input_c[0];
  assign cgp_core_016 = input_a[1] | input_c[1];
  assign cgp_core_017 = input_a[1] & input_c[1];
  assign cgp_core_018 = cgp_core_016 | cgp_core_015;
  assign cgp_core_019 = cgp_core_016 & input_a[0];
  assign cgp_core_020 = cgp_core_017 | cgp_core_019;
  assign cgp_core_021 = input_e[0] | input_f[0];
  assign cgp_core_022 = input_e[0] & input_f[0];
  assign cgp_core_023 = ~input_d[0];
  assign cgp_core_024 = input_a[1] ^ input_f[1];
  assign cgp_core_025 = input_f[1] | cgp_core_022;
  assign cgp_core_026 = input_f[1] & input_f[0];
  assign cgp_core_027 = input_e[1] | cgp_core_026;
  assign cgp_core_028 = input_b[0] & input_e[0];
  assign cgp_core_029 = input_d[0] & cgp_core_021;
  assign cgp_core_030 = input_d[1] | cgp_core_025;
  assign cgp_core_031 = input_d[1] & cgp_core_025;
  assign cgp_core_032 = cgp_core_030 | cgp_core_029;
  assign cgp_core_033 = cgp_core_030 & input_d[0];
  assign cgp_core_034 = cgp_core_031 | cgp_core_033;
  assign cgp_core_037 = ~(input_a[0] ^ input_c[1]);
  assign cgp_core_039 = cgp_core_018 | cgp_core_032;
  assign cgp_core_040 = cgp_core_018 & cgp_core_032;
  assign cgp_core_042 = cgp_core_039 & cgp_core_014;
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;
  assign cgp_core_044 = cgp_core_020 | cgp_core_034;
  assign cgp_core_046 = cgp_core_044 | cgp_core_043;
  assign cgp_core_047 = ~(input_e[0] & input_e[1]);
  assign cgp_core_048 = input_f[0] | input_b[1];
  assign cgp_core_051 = input_a[1] | input_b[1];
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_064 = input_b[1] & cgp_core_063;
  assign cgp_core_065 = cgp_core_064 & cgp_core_039;
  assign cgp_core_067 = input_d[1] ^ input_f[1];
  assign cgp_core_068 = cgp_core_058 | cgp_core_046;
  assign cgp_core_069 = cgp_core_065 | cgp_core_068;
  assign cgp_core_070 = ~(input_e[0] ^ input_a[1]);
  assign cgp_core_072 = cgp_core_069 | cgp_core_027;

  assign cgp_out[0] = cgp_core_072;
endmodule