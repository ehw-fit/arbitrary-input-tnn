module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070_not;
  wire cgp_core_071;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = ~(input_c[0] ^ input_a[1]);
  assign cgp_core_017 = ~(input_c[0] & input_b[1]);
  assign cgp_core_018 = input_f[1] | input_g[0];
  assign cgp_core_022 = ~(input_f[1] | input_f[0]);
  assign cgp_core_023 = input_d[1] ^ input_g[1];
  assign cgp_core_027 = input_b[0] ^ cgp_core_016;
  assign cgp_core_028 = input_b[0] ^ cgp_core_016;
  assign cgp_core_029 = input_d[1] | cgp_core_028;
  assign cgp_core_030 = cgp_core_022 ^ input_a[1];
  assign cgp_core_032 = ~(input_f[0] & input_c[0]);
  assign cgp_core_036 = ~(input_g[1] | input_a[0]);
  assign cgp_core_037 = ~input_c[1];
  assign cgp_core_038 = ~input_d[0];
  assign cgp_core_039 = input_e[0] ^ input_g[0];
  assign cgp_core_040 = ~(input_e[1] ^ input_f[1]);
  assign cgp_core_042 = ~(input_f[1] | input_d[0]);
  assign cgp_core_043 = input_e[1] & input_e[1];
  assign cgp_core_045 = input_a[1] | input_g[1];
  assign cgp_core_046 = input_c[0] ^ input_g[0];
  assign cgp_core_047 = cgp_core_032 ^ input_b[0];
  assign cgp_core_049 = ~(input_g[1] ^ input_b[1]);
  assign cgp_core_050_not = ~input_e[0];
  assign cgp_core_051 = input_d[0] & cgp_core_047;
  assign cgp_core_052 = cgp_core_049 ^ input_d[0];
  assign cgp_core_054 = ~(input_b[0] ^ cgp_core_045);
  assign cgp_core_055 = ~(input_f[1] & input_g[1]);
  assign cgp_core_056 = ~(input_e[0] & cgp_core_052);
  assign cgp_core_058 = input_e[0] & input_g[0];
  assign cgp_core_059 = ~(input_a[0] | cgp_core_058);
  assign cgp_core_061 = ~input_e[1];
  assign cgp_core_062 = input_d[1] & cgp_core_061;
  assign cgp_core_063 = input_f[1] & input_f[1];
  assign cgp_core_064 = ~(input_a[1] ^ input_a[0]);
  assign cgp_core_066 = input_b[0] & cgp_core_050_not;
  assign cgp_core_068 = ~input_c[0];
  assign cgp_core_069 = ~(cgp_core_027 ^ input_d[0]);
  assign cgp_core_070_not = ~input_g[1];
  assign cgp_core_071 = ~input_b[0];
  assign cgp_core_077 = cgp_core_059 | input_b[1];
  assign cgp_core_078 = input_e[1] ^ input_c[0];
  assign cgp_core_079 = input_a[0] | cgp_core_078;

  assign cgp_out[0] = 1'b0;
endmodule