module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_020_not;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046_not;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = input_d[0] ^ input_e[1];
  assign cgp_core_017 = input_d[0] & input_e[0];
  assign cgp_core_020_not = ~input_e[1];
  assign cgp_core_022_not = ~cgp_core_017;
  assign cgp_core_023 = input_e[1] ^ input_e[1];
  assign cgp_core_024 = input_a[0] & input_e[0];
  assign cgp_core_025 = input_a[1] ^ cgp_core_020_not;
  assign cgp_core_026_not = ~input_a[1];
  assign cgp_core_027 = ~(cgp_core_025 ^ cgp_core_024);
  assign cgp_core_028 = cgp_core_025 & cgp_core_024;
  assign cgp_core_030 = input_c[0] ^ input_g[0];
  assign cgp_core_031 = cgp_core_022_not & input_f[1];
  assign cgp_core_033 = input_b[0] & input_c[0];
  assign cgp_core_034 = input_b[1] ^ input_e[0];
  assign cgp_core_035 = ~(input_e[0] | input_g[1]);
  assign cgp_core_036 = input_e[0] ^ input_b[1];
  assign cgp_core_037 = input_d[0] ^ cgp_core_033;
  assign cgp_core_039 = ~(input_f[0] | input_g[0]);
  assign cgp_core_040 = input_b[1] & input_f[0];
  assign cgp_core_041 = ~input_f[1];
  assign cgp_core_042 = input_b[0] & input_g[1];
  assign cgp_core_043 = cgp_core_041 ^ input_c[1];
  assign cgp_core_044 = ~(cgp_core_041 & cgp_core_040);
  assign cgp_core_046_not = ~input_g[1];
  assign cgp_core_047 = input_c[1] & input_f[1];
  assign cgp_core_048 = input_c[1] ^ cgp_core_043;
  assign cgp_core_049 = input_g[0] & cgp_core_043;
  assign cgp_core_052 = ~(cgp_core_049 | input_d[0]);
  assign cgp_core_053 = input_c[0] ^ input_c[1];
  assign cgp_core_055 = cgp_core_053 ^ input_f[1];
  assign cgp_core_059 = cgp_core_031 | input_g[1];
  assign cgp_core_061 = ~(cgp_core_055 | input_g[0]);
  assign cgp_core_063 = cgp_core_030 & input_b[0];
  assign cgp_core_064 = ~(cgp_core_030 ^ input_e[1]);
  assign cgp_core_065 = ~(cgp_core_064 | input_g[0]);
  assign cgp_core_066 = cgp_core_048 & input_g[1];
  assign cgp_core_069 = ~(input_b[0] ^ cgp_core_048);
  assign cgp_core_070 = cgp_core_069 & cgp_core_065;
  assign cgp_core_071 = cgp_core_046_not | input_g[1];
  assign cgp_core_072 = input_d[0] & cgp_core_071;
  assign cgp_core_073 = ~(input_c[0] | cgp_core_070);
  assign cgp_core_074_not = ~input_d[0];
  assign cgp_core_075 = cgp_core_074_not & input_c[0];
  assign cgp_core_078 = ~cgp_core_063;
  assign cgp_core_079 = input_b[1] | input_g[1];

  assign cgp_out[0] = input_e[0];
endmodule