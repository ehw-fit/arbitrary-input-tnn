module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_045_not;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_096;

  assign cgp_core_018 = input_b[1] & input_f[1];
  assign cgp_core_019 = input_a[1] ^ input_e[1];
  assign cgp_core_022 = ~(input_f[1] ^ input_b[1]);
  assign cgp_core_023 = input_f[1] | input_b[1];
  assign cgp_core_024_not = ~input_a[0];
  assign cgp_core_025 = input_a[1] | input_g[0];
  assign cgp_core_027 = input_e[0] & input_d[1];
  assign cgp_core_028 = input_b[1] & input_d[1];
  assign cgp_core_029 = ~(input_d[0] | input_b[0]);
  assign cgp_core_030 = ~(input_b[1] | input_b[0]);
  assign cgp_core_031 = ~(input_b[1] | input_f[1]);
  assign cgp_core_032 = ~input_a[0];
  assign cgp_core_033 = input_d[1] & input_a[1];
  assign cgp_core_034 = ~input_b[0];
  assign cgp_core_035 = ~(input_h[0] & input_a[1]);
  assign cgp_core_037 = input_b[0] | input_g[0];
  assign cgp_core_039 = ~input_e[0];
  assign cgp_core_040 = input_c[1] | input_b[1];
  assign cgp_core_041 = ~(input_b[0] & input_d[0]);
  assign cgp_core_045_not = ~input_b[1];
  assign cgp_core_046 = ~(input_f[1] ^ input_b[1]);
  assign cgp_core_047 = input_a[1] & input_f[1];
  assign cgp_core_048 = input_h[1] & input_a[1];
  assign cgp_core_049 = input_a[0] & input_d[1];
  assign cgp_core_052 = ~(input_a[0] | input_h[1]);
  assign cgp_core_054 = input_g[0] ^ input_e[0];
  assign cgp_core_055 = ~(input_h[0] | input_b[1]);
  assign cgp_core_056 = ~input_b[0];
  assign cgp_core_057 = ~(input_f[1] ^ input_f[1]);
  assign cgp_core_058 = ~(input_g[1] ^ input_e[0]);
  assign cgp_core_059 = ~(input_h[0] ^ input_h[1]);
  assign cgp_core_060 = ~(input_c[0] | input_d[1]);
  assign cgp_core_064 = cgp_core_040 | input_f[1];
  assign cgp_core_065 = input_c[1] & input_f[1];
  assign cgp_core_066 = cgp_core_064 | input_e[1];
  assign cgp_core_067 = input_b[1] & input_e[1];
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = input_g[1] | cgp_core_068;
  assign cgp_core_071 = input_e[0] | input_g[1];
  assign cgp_core_072 = input_c[1] ^ input_a[1];
  assign cgp_core_073 = ~cgp_core_069;
  assign cgp_core_074 = cgp_core_033 & cgp_core_073;
  assign cgp_core_076 = input_d[1] & input_b[1];
  assign cgp_core_077 = ~(input_a[0] | input_a[0]);
  assign cgp_core_078 = ~cgp_core_066;
  assign cgp_core_079 = input_h[1] & cgp_core_078;
  assign cgp_core_083 = ~input_a[0];
  assign cgp_core_085 = input_d[1] & input_d[1];
  assign cgp_core_087 = ~(input_h[0] & input_b[0]);
  assign cgp_core_088 = input_c[1] | input_g[1];
  assign cgp_core_091 = ~(input_h[0] | input_e[1]);
  assign cgp_core_092 = ~(input_g[0] & input_f[1]);
  assign cgp_core_096 = cgp_core_079 | cgp_core_074;

  assign cgp_out[0] = cgp_core_096;
endmodule