module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097_not;
  wire cgp_core_098;

  assign cgp_core_020 = ~(input_c[0] & input_e[0]);
  assign cgp_core_021 = input_c[0] & input_e[0];
  assign cgp_core_022 = ~(input_c[1] & input_e[1]);
  assign cgp_core_023 = input_c[1] & input_e[1];
  assign cgp_core_024 = ~cgp_core_022;
  assign cgp_core_025 = cgp_core_022 ^ cgp_core_021;
  assign cgp_core_026 = cgp_core_023 | input_d[2];
  assign cgp_core_027_not = ~input_c[2];
  assign cgp_core_029 = ~(input_f[2] ^ cgp_core_026);
  assign cgp_core_032 = input_e[2] ^ cgp_core_020;
  assign cgp_core_034 = input_d[1] ^ cgp_core_024;
  assign cgp_core_035 = input_a[2] & cgp_core_024;
  assign cgp_core_039 = input_a[0] & cgp_core_029;
  assign cgp_core_040 = input_a[2] & input_f[1];
  assign cgp_core_041_not = ~cgp_core_039;
  assign cgp_core_042 = cgp_core_039 & input_e[0];
  assign cgp_core_044 = input_f[1] ^ cgp_core_040;
  assign cgp_core_047 = input_d[0] & input_f[0];
  assign cgp_core_048 = input_c[0] | input_f[1];
  assign cgp_core_049 = input_d[1] & input_f[1];
  assign cgp_core_050 = cgp_core_048 ^ cgp_core_047;
  assign cgp_core_051 = cgp_core_048 & input_b[1];
  assign cgp_core_052 = input_a[2] & cgp_core_051;
  assign cgp_core_053 = input_d[0] ^ input_f[2];
  assign cgp_core_054 = input_e[1] & input_a[0];
  assign cgp_core_055 = ~(cgp_core_053 & cgp_core_052);
  assign cgp_core_056 = input_b[0] & cgp_core_052;
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_060 = ~(input_b[1] | cgp_core_050);
  assign cgp_core_061 = ~input_b[1];
  assign cgp_core_063 = cgp_core_060 & input_b[0];
  assign cgp_core_064 = cgp_core_061 | cgp_core_063;
  assign cgp_core_065 = input_b[2] & input_d[1];
  assign cgp_core_066 = input_b[2] & input_e[2];
  assign cgp_core_067 = cgp_core_065 ^ cgp_core_064;
  assign cgp_core_068 = cgp_core_065 & input_f[1];
  assign cgp_core_069 = input_e[0] & cgp_core_068;
  assign cgp_core_070 = cgp_core_057 ^ input_b[2];
  assign cgp_core_075 = ~(cgp_core_070 ^ input_f[2]);
  assign cgp_core_076 = cgp_core_044 & cgp_core_075;
  assign cgp_core_078 = ~(input_f[1] ^ cgp_core_070);
  assign cgp_core_080 = ~input_b[0];
  assign cgp_core_081 = input_a[1] & input_b[0];
  assign cgp_core_083 = ~(cgp_core_041_not ^ cgp_core_067);
  assign cgp_core_085 = ~input_c[0];
  assign cgp_core_086 = input_f[2] & cgp_core_085;
  assign cgp_core_087 = cgp_core_086 & input_c[1];
  assign cgp_core_088 = ~(input_d[0] ^ cgp_core_060);
  assign cgp_core_090 = ~input_a[2];
  assign cgp_core_091 = cgp_core_032 & input_f[0];
  assign cgp_core_093 = ~(cgp_core_032 ^ input_a[2]);
  assign cgp_core_095 = cgp_core_087 | cgp_core_081;
  assign cgp_core_096 = ~(input_d[0] ^ cgp_core_095);
  assign cgp_core_097_not = ~cgp_core_093;
  assign cgp_core_098 = input_b[2] | input_e[2];

  assign cgp_out[0] = 1'b1;
endmodule