module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_012 = input_b[0] ^ input_d[0];
  assign cgp_core_013 = input_b[0] & input_d[0];
  assign cgp_core_014 = input_b[1] ^ input_d[1];
  assign cgp_core_015 = input_b[1] & input_d[1];
  assign cgp_core_016 = cgp_core_014 ^ cgp_core_013;
  assign cgp_core_017 = cgp_core_014 & cgp_core_013;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = input_c[0] ^ input_e[0];
  assign cgp_core_020 = input_c[0] & input_e[0];
  assign cgp_core_021 = input_c[1] ^ input_e[1];
  assign cgp_core_022 = input_c[1] & input_e[1];
  assign cgp_core_023 = cgp_core_021 ^ cgp_core_020;
  assign cgp_core_024 = cgp_core_021 & cgp_core_020;
  assign cgp_core_025 = cgp_core_022 | cgp_core_024;
  assign cgp_core_027 = input_a[0] & cgp_core_019;
  assign cgp_core_028 = input_a[1] ^ cgp_core_023;
  assign cgp_core_029 = input_a[1] & cgp_core_023;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_033 = cgp_core_025 | cgp_core_032;
  assign cgp_core_034 = cgp_core_025 & input_a[1];
  assign cgp_core_035 = input_e[0] | input_e[0];
  assign cgp_core_036 = ~cgp_core_034;
  assign cgp_core_037 = ~cgp_core_033;
  assign cgp_core_038 = cgp_core_018 & cgp_core_037;
  assign cgp_core_040 = ~(cgp_core_018 ^ cgp_core_033);
  assign cgp_core_041 = cgp_core_040 & cgp_core_036;
  assign cgp_core_042 = ~cgp_core_030;
  assign cgp_core_043 = cgp_core_016 & cgp_core_042;
  assign cgp_core_044 = cgp_core_043 & cgp_core_041;
  assign cgp_core_045 = ~(cgp_core_016 ^ cgp_core_030);
  assign cgp_core_046 = cgp_core_045 & cgp_core_041;
  assign cgp_core_047 = input_b[0] | input_e[1];
  assign cgp_core_051 = cgp_core_012 & cgp_core_046;
  assign cgp_core_053 = cgp_core_038 | cgp_core_051;
  assign cgp_core_054 = cgp_core_044 | cgp_core_053;

  assign cgp_out[0] = cgp_core_054;
endmodule