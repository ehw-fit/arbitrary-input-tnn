module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033_not;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;

  assign cgp_core_017 = input_b[0] ^ input_c[0];
  assign cgp_core_018 = input_a[1] & input_c[0];
  assign cgp_core_019_not = ~input_b[1];
  assign cgp_core_020 = input_b[1] & input_b[2];
  assign cgp_core_021 = ~(input_e[2] ^ cgp_core_018);
  assign cgp_core_022 = ~(input_b[2] ^ input_d[0]);
  assign cgp_core_023 = ~input_c[1];
  assign cgp_core_024 = input_b[2] ^ input_c[2];
  assign cgp_core_025 = input_a[0] & input_b[2];
  assign cgp_core_026 = ~(input_e[1] & input_b[1]);
  assign cgp_core_027 = cgp_core_024 & input_d[1];
  assign cgp_core_029 = input_d[0] ^ input_e[0];
  assign cgp_core_031 = ~(input_d[1] ^ input_e[1]);
  assign cgp_core_033_not = ~cgp_core_031;
  assign cgp_core_035 = input_d[1] | input_c[0];
  assign cgp_core_036 = ~(input_d[2] & input_c[1]);
  assign cgp_core_037 = ~(input_d[2] ^ input_e[2]);
  assign cgp_core_038 = input_c[0] ^ cgp_core_035;
  assign cgp_core_039 = cgp_core_036 & cgp_core_035;
  assign cgp_core_041 = cgp_core_017 ^ cgp_core_029;
  assign cgp_core_042 = ~(cgp_core_017 | input_d[1]);
  assign cgp_core_043 = ~(cgp_core_021 | input_b[2]);
  assign cgp_core_044 = input_d[2] & cgp_core_033_not;
  assign cgp_core_045 = input_b[0] ^ input_d[2];
  assign cgp_core_046 = input_e[1] & cgp_core_042;
  assign cgp_core_047 = ~cgp_core_044;
  assign cgp_core_048 = cgp_core_026 ^ input_b[2];
  assign cgp_core_049 = ~input_a[0];
  assign cgp_core_050 = input_b[2] ^ input_d[2];
  assign cgp_core_051 = cgp_core_048 & cgp_core_047;
  assign cgp_core_052 = cgp_core_049 & cgp_core_051;
  assign cgp_core_053 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_054 = ~(input_b[0] & input_d[0]);
  assign cgp_core_056 = cgp_core_053 & cgp_core_052;
  assign cgp_core_057 = ~(cgp_core_054 | cgp_core_056);
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_063 = ~input_c[2];
  assign cgp_core_064 = input_a[2] & cgp_core_063;
  assign cgp_core_066 = input_a[2] | cgp_core_050;
  assign cgp_core_068 = ~cgp_core_045;
  assign cgp_core_069 = input_a[1] & cgp_core_068;
  assign cgp_core_070 = cgp_core_069 & input_c[1];
  assign cgp_core_071 = input_a[1] & cgp_core_045;
  assign cgp_core_073 = ~input_d[0];
  assign cgp_core_074 = input_a[0] & cgp_core_073;
  assign cgp_core_075 = input_a[0] & input_b[0];
  assign cgp_core_076 = ~(input_a[0] ^ input_d[0]);

  assign cgp_out[0] = 1'b0;
endmodule