module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060_not;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079_not;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_097;
  wire cgp_core_099;

  assign cgp_core_020 = ~(input_b[2] ^ input_f[2]);
  assign cgp_core_024 = input_e[0] ^ input_f[2];
  assign cgp_core_025_not = ~input_d[2];
  assign cgp_core_026 = ~(input_e[0] ^ input_a[2]);
  assign cgp_core_027 = ~input_a[0];
  assign cgp_core_028 = input_b[2] & input_b[2];
  assign cgp_core_030 = input_b[2] ^ input_a[2];
  assign cgp_core_031 = input_d[0] & input_b[2];
  assign cgp_core_032 = input_b[0] | input_c[2];
  assign cgp_core_033 = input_f[1] | input_a[2];
  assign cgp_core_037 = ~input_b[0];
  assign cgp_core_038 = input_b[1] | input_c[0];
  assign cgp_core_039 = ~input_b[0];
  assign cgp_core_040_not = ~input_f[0];
  assign cgp_core_041 = ~input_e[0];
  assign cgp_core_042 = input_d[0] & input_a[2];
  assign cgp_core_044 = ~input_f[1];
  assign cgp_core_045 = input_c[2] ^ input_c[0];
  assign cgp_core_047 = ~(input_f[2] ^ input_e[0]);
  assign cgp_core_051 = ~(input_f[1] ^ input_e[0]);
  assign cgp_core_053 = ~(input_d[2] ^ input_c[1]);
  assign cgp_core_054 = ~(input_d[2] & input_e[0]);
  assign cgp_core_055 = input_e[0] & input_c[0];
  assign cgp_core_056 = input_d[2] ^ input_f[2];
  assign cgp_core_057 = ~(input_d[0] | input_b[2]);
  assign cgp_core_060_not = ~input_d[1];
  assign cgp_core_061 = input_e[1] & input_e[2];
  assign cgp_core_062 = input_a[1] & input_a[1];
  assign cgp_core_064 = ~(input_e[1] ^ input_b[2]);
  assign cgp_core_065 = input_d[2] ^ input_a[1];
  assign cgp_core_066 = input_b[0] & input_a[1];
  assign cgp_core_067 = input_e[1] | input_b[2];
  assign cgp_core_068 = ~(input_d[0] | input_a[2]);
  assign cgp_core_069 = input_a[2] | input_b[1];
  assign cgp_core_070 = ~input_c[2];
  assign cgp_core_071 = ~(input_b[2] | input_a[2]);
  assign cgp_core_072 = ~(input_b[1] ^ input_f[2]);
  assign cgp_core_074 = ~(input_d[2] ^ input_e[0]);
  assign cgp_core_075 = ~(input_b[2] ^ input_c[0]);
  assign cgp_core_076 = input_a[2] & input_e[2];
  assign cgp_core_078 = ~(input_d[1] | input_c[2]);
  assign cgp_core_079_not = ~input_e[2];
  assign cgp_core_080 = ~input_b[2];
  assign cgp_core_081 = ~(input_f[2] & input_f[0]);
  assign cgp_core_082 = ~input_d[0];
  assign cgp_core_083 = input_a[0] | input_d[1];
  assign cgp_core_084 = ~(input_c[2] | input_d[2]);
  assign cgp_core_085 = input_c[0] & input_f[1];
  assign cgp_core_086 = ~(input_d[1] ^ input_d[2]);
  assign cgp_core_088 = ~input_d[1];
  assign cgp_core_089 = ~input_d[2];
  assign cgp_core_091 = ~(input_d[2] ^ input_d[2]);
  assign cgp_core_092 = ~(input_e[2] ^ input_d[1]);
  assign cgp_core_093 = ~(input_e[0] ^ input_f[0]);
  assign cgp_core_094 = ~input_f[1];
  assign cgp_core_097 = ~(input_d[2] & input_b[0]);
  assign cgp_core_099 = input_c[2] | cgp_core_076;

  assign cgp_out[0] = cgp_core_099;
endmodule