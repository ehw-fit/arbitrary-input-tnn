module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_048_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_054_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061_not;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_014 = ~(input_c[1] & input_a[1]);
  assign cgp_core_018 = ~(input_b[0] ^ input_e[1]);
  assign cgp_core_019 = input_d[0] & input_f[1];
  assign cgp_core_020 = ~(input_f[1] | input_a[0]);
  assign cgp_core_021 = ~(input_e[0] ^ input_b[0]);
  assign cgp_core_023_not = ~input_e[1];
  assign cgp_core_024 = ~input_d[1];
  assign cgp_core_025 = ~(input_a[1] | input_d[0]);
  assign cgp_core_026 = input_e[1] ^ input_e[0];
  assign cgp_core_027 = input_a[0] ^ input_f[1];
  assign cgp_core_030 = ~input_e[0];
  assign cgp_core_032_not = ~input_b[0];
  assign cgp_core_033 = ~(input_c[1] ^ input_d[1]);
  assign cgp_core_035 = ~(input_f[1] ^ input_a[1]);
  assign cgp_core_036_not = ~input_c[0];
  assign cgp_core_040 = ~(input_b[1] & input_e[1]);
  assign cgp_core_041 = input_e[1] | input_e[1];
  assign cgp_core_042 = ~input_d[1];
  assign cgp_core_043 = input_c[0] | input_f[0];
  assign cgp_core_046 = input_e[1] | cgp_core_043;
  assign cgp_core_048_not = ~input_a[0];
  assign cgp_core_049 = input_a[0] & input_c[1];
  assign cgp_core_050 = ~(input_f[1] & input_e[0]);
  assign cgp_core_051 = ~(input_f[1] ^ input_a[0]);
  assign cgp_core_054_not = ~input_e[1];
  assign cgp_core_056 = input_c[0] | input_e[1];
  assign cgp_core_057 = input_e[0] | input_c[0];
  assign cgp_core_058 = ~input_d[1];
  assign cgp_core_061_not = ~input_c[0];
  assign cgp_core_062 = ~(input_d[0] | input_c[0]);
  assign cgp_core_064 = ~(input_b[0] & input_a[0]);
  assign cgp_core_068 = input_a[1] | cgp_core_046;
  assign cgp_core_069 = input_c[1] | cgp_core_068;
  assign cgp_core_070 = input_d[1] | input_e[0];
  assign cgp_core_071 = input_f[1] | cgp_core_070;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;

  assign cgp_out[0] = cgp_core_072;
endmodule