module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061_not;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_081;
  wire cgp_core_082_not;

  assign cgp_core_016 = input_a[0] | input_g[1];
  assign cgp_core_017 = input_a[0] | input_d[0];
  assign cgp_core_018 = ~input_c[0];
  assign cgp_core_020 = input_c[0] ^ input_b[0];
  assign cgp_core_021 = input_e[1] & input_e[1];
  assign cgp_core_022 = ~(input_f[0] | cgp_core_021);
  assign cgp_core_023 = input_e[0] ^ input_f[1];
  assign cgp_core_025 = ~input_a[1];
  assign cgp_core_026 = input_c[0] & input_c[1];
  assign cgp_core_030 = ~(input_d[0] | input_e[1]);
  assign cgp_core_031 = ~(input_a[0] ^ input_a[1]);
  assign cgp_core_034 = input_e[0] ^ cgp_core_031;
  assign cgp_core_035 = input_f[1] & cgp_core_031;
  assign cgp_core_038 = cgp_core_026 & input_f[0];
  assign cgp_core_039 = cgp_core_016 ^ input_f[0];
  assign cgp_core_040 = ~(input_b[0] | cgp_core_030);
  assign cgp_core_041 = ~(cgp_core_020 & input_e[1]);
  assign cgp_core_042 = ~(input_c[1] & cgp_core_034);
  assign cgp_core_043 = ~(input_b[0] & cgp_core_040);
  assign cgp_core_044 = ~(input_b[0] ^ input_a[1]);
  assign cgp_core_045 = ~(cgp_core_042 ^ cgp_core_044);
  assign cgp_core_046 = input_d[1] ^ input_f[0];
  assign cgp_core_047 = input_c[1] | input_e[0];
  assign cgp_core_048 = ~cgp_core_046;
  assign cgp_core_053 = ~(input_b[0] ^ input_f[0]);
  assign cgp_core_054 = input_b[0] & input_f[0];
  assign cgp_core_055 = ~(input_a[1] | input_e[0]);
  assign cgp_core_058 = ~(input_e[0] ^ cgp_core_054);
  assign cgp_core_059 = input_c[1] | input_g[0];
  assign cgp_core_061_not = ~input_c[1];
  assign cgp_core_062 = ~input_c[0];
  assign cgp_core_063 = cgp_core_062 & input_b[1];
  assign cgp_core_064 = ~(cgp_core_059 ^ input_c[0]);
  assign cgp_core_065 = input_g[1] | cgp_core_064;
  assign cgp_core_066 = cgp_core_065 & input_a[0];
  assign cgp_core_067 = ~(input_f[0] ^ cgp_core_059);
  assign cgp_core_068 = cgp_core_067 & input_b[0];
  assign cgp_core_070 = cgp_core_043 & input_b[1];
  assign cgp_core_071 = input_g[1] & input_a[0];
  assign cgp_core_073 = cgp_core_043 & input_a[0];
  assign cgp_core_075 = input_g[1] & input_b[0];
  assign cgp_core_076 = cgp_core_075 ^ input_g[1];
  assign cgp_core_077 = ~(cgp_core_039 ^ cgp_core_053);
  assign cgp_core_081 = ~(input_b[0] & input_c[0]);
  assign cgp_core_082_not = ~cgp_core_061_not;

  assign cgp_out[0] = 1'b1;
endmodule