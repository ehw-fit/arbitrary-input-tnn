module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;

  assign cgp_core_018 = input_d[1] | input_e[1];
  assign cgp_core_019 = input_d[1] & input_e[1];
  assign cgp_core_021 = cgp_core_018 & input_e[0];
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_027 = input_g[0] ^ input_d[1];
  assign cgp_core_028 = input_d[1] & input_g[0];
  assign cgp_core_029 = input_g[1] & input_b[0];
  assign cgp_core_030 = cgp_core_022 | input_a[1];
  assign cgp_core_031 = cgp_core_022 & input_a[1];
  assign cgp_core_032 = input_d[1] | input_e[1];
  assign cgp_core_033 = ~(input_a[1] & input_c[1]);
  assign cgp_core_034 = ~input_g[0];
  assign cgp_core_036 = input_d[1] ^ input_c[1];
  assign cgp_core_037 = ~(input_g[0] ^ input_g[0]);
  assign cgp_core_038 = input_g[0] ^ input_g[1];
  assign cgp_core_044 = ~(input_b[1] | input_d[0]);
  assign cgp_core_045 = input_g[0] | input_a[1];
  assign cgp_core_047 = input_g[1] | input_f[1];
  assign cgp_core_048 = input_f[1] & input_a[1];
  assign cgp_core_049 = input_g[0] ^ input_d[1];
  assign cgp_core_050_not = ~input_c[0];
  assign cgp_core_052 = input_g[1] | input_f[1];
  assign cgp_core_053 = ~(input_b[0] | input_f[0]);
  assign cgp_core_054 = input_g[1] & input_f[1];
  assign cgp_core_056 = input_b[1] & cgp_core_052;
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = cgp_core_031 & cgp_core_058;
  assign cgp_core_060 = ~(input_c[1] | cgp_core_057);
  assign cgp_core_063 = cgp_core_030 & cgp_core_060;
  assign cgp_core_064 = ~(input_f[0] & input_f[0]);
  assign cgp_core_065 = ~(input_d[1] | input_b[1]);
  assign cgp_core_067 = ~(input_c[1] | input_g[0]);
  assign cgp_core_068 = input_a[0] | input_g[1];
  assign cgp_core_070 = ~(input_a[0] & input_g[1]);
  assign cgp_core_072 = input_e[0] & input_b[0];
  assign cgp_core_073 = ~(input_c[0] ^ input_c[0]);
  assign cgp_core_074 = input_e[0] | input_b[0];
  assign cgp_core_075 = input_c[1] | input_e[1];
  assign cgp_core_076 = ~(input_b[1] | input_b[1]);
  assign cgp_core_078 = cgp_core_063 | cgp_core_059;

  assign cgp_out[0] = cgp_core_078;
endmodule