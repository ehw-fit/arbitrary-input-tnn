module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067_not;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071_not;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_092;
  wire cgp_core_094;
  wire cgp_core_095;

  assign cgp_core_018 = input_b[0] ^ input_c[0];
  assign cgp_core_019 = ~(input_h[1] | input_c[0]);
  assign cgp_core_021 = input_g[0] & input_c[1];
  assign cgp_core_022 = ~(input_h[0] & cgp_core_019);
  assign cgp_core_025 = ~(input_a[0] & cgp_core_018);
  assign cgp_core_027 = input_b[1] ^ cgp_core_022;
  assign cgp_core_028 = input_a[1] & cgp_core_022;
  assign cgp_core_032 = input_c[0] ^ input_e[1];
  assign cgp_core_034 = input_g[0] ^ input_h[0];
  assign cgp_core_035 = ~(input_g[0] & input_d[0]);
  assign cgp_core_036 = ~(input_g[1] | input_a[0]);
  assign cgp_core_037 = input_g[1] & input_h[1];
  assign cgp_core_038 = input_e[0] ^ cgp_core_035;
  assign cgp_core_039 = input_a[1] & cgp_core_035;
  assign cgp_core_040 = input_b[0] | cgp_core_039;
  assign cgp_core_043 = input_d[1] ^ input_d[1];
  assign cgp_core_044 = input_d[1] & input_g[0];
  assign cgp_core_046 = cgp_core_043 & cgp_core_034;
  assign cgp_core_048 = cgp_core_040 ^ cgp_core_044;
  assign cgp_core_049 = cgp_core_040 & input_f[1];
  assign cgp_core_051 = cgp_core_025 & input_c[1];
  assign cgp_core_053 = ~(input_b[1] | input_g[0]);
  assign cgp_core_055 = cgp_core_027 | input_d[0];
  assign cgp_core_057 = ~(cgp_core_032 ^ cgp_core_048);
  assign cgp_core_061 = ~(input_b[0] | input_e[0]);
  assign cgp_core_063 = input_f[0] & input_g[0];
  assign cgp_core_064 = input_c[1] ^ cgp_core_061;
  assign cgp_core_065 = input_c[1] & input_c[1];
  assign cgp_core_066 = input_c[1] | input_d[1];
  assign cgp_core_067_not = ~input_f[0];
  assign cgp_core_069 = input_e[1] | input_f[1];
  assign cgp_core_070 = input_e[1] & input_f[1];
  assign cgp_core_071_not = ~input_h[1];
  assign cgp_core_072 = ~(cgp_core_069 | input_h[0]);
  assign cgp_core_073 = cgp_core_070 | input_a[0];
  assign cgp_core_078 = ~cgp_core_073;
  assign cgp_core_079 = input_g[0] & cgp_core_078;
  assign cgp_core_081 = ~(cgp_core_057 ^ cgp_core_073);
  assign cgp_core_083 = ~cgp_core_071_not;
  assign cgp_core_084 = cgp_core_051 & input_f[1];
  assign cgp_core_086 = ~(input_f[1] ^ cgp_core_071_not);
  assign cgp_core_087 = input_a[1] & input_e[1];
  assign cgp_core_092 = ~(input_f[1] | cgp_core_087);
  assign cgp_core_094 = cgp_core_087 | input_b[1];
  assign cgp_core_095 = cgp_core_066 | input_a[0];

  assign cgp_out[0] = 1'b1;
endmodule