module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_082;
  wire cgp_core_083;

  assign cgp_core_016 = ~(input_b[1] | input_a[1]);
  assign cgp_core_017 = ~input_c[1];
  assign cgp_core_018 = input_a[1] | input_c[1];
  assign cgp_core_019 = input_a[1] & input_c[1];
  assign cgp_core_020 = cgp_core_018 | input_d[0];
  assign cgp_core_021 = input_c[0] & input_a[0];
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_024_not = ~input_g[1];
  assign cgp_core_025 = input_e[1] | input_g[1];
  assign cgp_core_026 = input_e[1] & input_g[1];
  assign cgp_core_028 = cgp_core_025 & input_e[0];
  assign cgp_core_029 = cgp_core_026 | cgp_core_028;
  assign cgp_core_030 = ~(input_f[0] & input_a[1]);
  assign cgp_core_033 = input_d[1] & cgp_core_025;
  assign cgp_core_034 = input_d[0] | input_d[1];
  assign cgp_core_035 = input_g[0] | input_g[0];
  assign cgp_core_037 = cgp_core_029 | cgp_core_033;
  assign cgp_core_038 = input_e[0] & input_d[1];
  assign cgp_core_039 = ~input_g[1];
  assign cgp_core_041 = ~cgp_core_020;
  assign cgp_core_044 = ~cgp_core_041;
  assign cgp_core_045 = input_g[0] | cgp_core_044;
  assign cgp_core_048 = input_a[0] | cgp_core_045;
  assign cgp_core_049 = cgp_core_022 & cgp_core_045;
  assign cgp_core_050 = cgp_core_037 | cgp_core_049;
  assign cgp_core_053 = ~(input_c[0] ^ input_b[0]);
  assign cgp_core_055 = input_g[1] ^ input_e[0];
  assign cgp_core_056 = input_b[1] & input_f[1];
  assign cgp_core_058 = ~(input_c[1] & input_g[1]);
  assign cgp_core_060 = ~(input_f[0] | input_d[1]);
  assign cgp_core_062 = input_b[0] | input_f[1];
  assign cgp_core_063 = input_e[0] ^ input_d[0];
  assign cgp_core_064 = ~cgp_core_056;
  assign cgp_core_065 = cgp_core_048 & cgp_core_064;
  assign cgp_core_067 = ~(input_d[1] | input_f[1]);
  assign cgp_core_068 = input_d[0] ^ input_g[1];
  assign cgp_core_069_not = ~input_f[1];
  assign cgp_core_074 = ~(input_a[0] ^ input_e[0]);
  assign cgp_core_075 = ~input_c[0];
  assign cgp_core_077 = input_c[0] ^ input_d[1];
  assign cgp_core_078 = input_d[1] & input_f[1];
  assign cgp_core_082 = cgp_core_050 | cgp_core_038;
  assign cgp_core_083 = cgp_core_065 | cgp_core_082;

  assign cgp_out[0] = cgp_core_083;
endmodule