module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062_not;
  wire cgp_core_063;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_080;

  assign cgp_core_017 = ~(input_d[2] ^ input_d[2]);
  assign cgp_core_018 = input_d[2] ^ input_d[1];
  assign cgp_core_020 = ~(input_e[0] | input_a[0]);
  assign cgp_core_021 = ~input_b[1];
  assign cgp_core_023 = input_b[1] | input_a[1];
  assign cgp_core_024 = input_a[2] | input_b[2];
  assign cgp_core_025 = input_a[2] & input_b[2];
  assign cgp_core_027 = cgp_core_024 & cgp_core_023;
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_029 = ~(input_d[2] & input_b[1]);
  assign cgp_core_032 = input_a[2] ^ input_a[0];
  assign cgp_core_033 = ~(input_e[2] ^ input_e[0]);
  assign cgp_core_034 = input_b[0] & input_d[0];
  assign cgp_core_036 = input_e[1] & input_a[2];
  assign cgp_core_037 = input_c[1] & input_a[1];
  assign cgp_core_039 = ~(input_e[2] ^ input_e[2]);
  assign cgp_core_040 = input_d[2] | input_e[2];
  assign cgp_core_043 = ~input_c[2];
  assign cgp_core_044 = ~(input_d[2] ^ input_a[2]);
  assign cgp_core_045 = ~(input_d[2] & input_d[0]);
  assign cgp_core_046 = input_c[0] ^ input_e[0];
  assign cgp_core_047 = ~(input_a[2] ^ input_b[2]);
  assign cgp_core_050 = input_c[2] | input_c[0];
  assign cgp_core_052 = ~(input_b[0] ^ input_a[1]);
  assign cgp_core_054 = cgp_core_040 & input_c[2];
  assign cgp_core_055 = input_c[2] & input_c[1];
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_057 = input_a[1] | input_d[2];
  assign cgp_core_058 = ~(input_e[1] ^ input_b[2]);
  assign cgp_core_059 = ~input_d[2];
  assign cgp_core_061 = cgp_core_028 & cgp_core_056;
  assign cgp_core_062_not = ~input_c[2];
  assign cgp_core_063 = ~(input_c[0] | input_c[0]);
  assign cgp_core_067 = ~input_e[2];
  assign cgp_core_069 = ~(input_d[1] ^ input_d[2]);
  assign cgp_core_070 = ~(input_d[2] & input_e[2]);
  assign cgp_core_071 = cgp_core_070 & cgp_core_061;
  assign cgp_core_073 = input_b[2] ^ input_e[0];
  assign cgp_core_076 = ~input_c[1];
  assign cgp_core_077 = ~(input_b[2] & input_d[1]);
  assign cgp_core_080 = ~(input_c[1] | input_a[0]);

  assign cgp_out[0] = cgp_core_071;
endmodule