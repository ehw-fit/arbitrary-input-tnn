module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056_not;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077_not;

  assign cgp_core_016 = input_a[0] ^ input_d[0];
  assign cgp_core_017 = ~(input_b[1] & input_e[1]);
  assign cgp_core_018 = input_c[0] & input_d[1];
  assign cgp_core_020 = cgp_core_018 | input_b[1];
  assign cgp_core_023 = input_e[1] ^ input_g[0];
  assign cgp_core_029 = ~(input_d[1] & input_g[0]);
  assign cgp_core_030 = ~cgp_core_016;
  assign cgp_core_031 = ~(cgp_core_016 & cgp_core_023);
  assign cgp_core_032 = ~(input_f[1] | input_d[0]);
  assign cgp_core_033 = input_g[1] & input_b[0];
  assign cgp_core_034 = ~(cgp_core_032 ^ input_e[1]);
  assign cgp_core_035 = ~(input_d[0] | cgp_core_031);
  assign cgp_core_036 = input_g[0] | cgp_core_035;
  assign cgp_core_037 = ~(input_e[1] & input_a[0]);
  assign cgp_core_038 = ~(input_b[0] & cgp_core_029);
  assign cgp_core_039 = ~(input_g[0] ^ input_b[1]);
  assign cgp_core_040 = cgp_core_037 & input_c[0];
  assign cgp_core_041 = input_a[0] | input_b[1];
  assign cgp_core_042 = ~input_g[0];
  assign cgp_core_043 = input_g[0] & input_c[0];
  assign cgp_core_044 = input_f[1] | input_g[0];
  assign cgp_core_046 = input_b[0] ^ input_g[1];
  assign cgp_core_047 = ~(cgp_core_044 ^ cgp_core_043);
  assign cgp_core_049 = input_a[0] | input_d[1];
  assign cgp_core_050 = input_g[0] & input_b[1];
  assign cgp_core_051 = ~(input_a[1] ^ input_c[0]);
  assign cgp_core_052 = ~(input_a[1] | input_b[1]);
  assign cgp_core_053 = input_e[1] ^ input_c[1];
  assign cgp_core_054 = ~input_f[0];
  assign cgp_core_056_not = ~input_b[1];
  assign cgp_core_058 = input_b[0] & input_e[0];
  assign cgp_core_059 = input_d[1] & input_f[0];
  assign cgp_core_060 = input_d[0] & input_f[1];
  assign cgp_core_061 = input_b[0] | input_a[1];
  assign cgp_core_063 = ~input_a[0];
  assign cgp_core_064 = input_e[1] & input_g[0];
  assign cgp_core_066 = ~cgp_core_053;
  assign cgp_core_069 = input_a[0] | input_d[1];
  assign cgp_core_070 = ~(input_a[0] & cgp_core_064);
  assign cgp_core_071 = ~(input_c[0] & input_e[1]);
  assign cgp_core_072 = ~input_e[1];
  assign cgp_core_074 = ~cgp_core_030;
  assign cgp_core_075 = cgp_core_074 | input_f[0];
  assign cgp_core_077_not = ~cgp_core_059;

  assign cgp_out[0] = input_b[0];
endmodule