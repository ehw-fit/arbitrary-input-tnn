module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_057_not;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;

  assign cgp_core_016 = input_f[1] ^ input_g[0];
  assign cgp_core_017 = input_d[1] & input_f[0];
  assign cgp_core_019 = input_a[0] | input_e[1];
  assign cgp_core_020 = input_c[0] & input_b[1];
  assign cgp_core_021 = ~(input_g[1] & input_b[0]);
  assign cgp_core_022 = input_d[1] & input_d[1];
  assign cgp_core_023 = input_e[1] ^ input_c[1];
  assign cgp_core_024 = input_g[0] | input_e[1];
  assign cgp_core_025 = input_d[1] ^ input_g[1];
  assign cgp_core_028 = ~(input_c[1] ^ input_d[1]);
  assign cgp_core_029 = input_b[0] ^ input_e[0];
  assign cgp_core_030 = ~(input_f[0] & cgp_core_023);
  assign cgp_core_032 = ~(input_d[1] & input_f[1]);
  assign cgp_core_033 = ~input_c[0];
  assign cgp_core_034 = ~(input_f[1] & input_d[0]);
  assign cgp_core_035_not = ~input_f[1];
  assign cgp_core_037 = ~(cgp_core_029 | input_c[1]);
  assign cgp_core_038 = ~input_b[1];
  assign cgp_core_042 = input_c[0] ^ input_d[0];
  assign cgp_core_043_not = ~input_a[0];
  assign cgp_core_044 = input_a[0] & input_f[0];
  assign cgp_core_046 = ~(input_c[1] & input_g[1]);
  assign cgp_core_047 = input_f[1] & input_d[1];
  assign cgp_core_051 = cgp_core_038 ^ input_g[0];
  assign cgp_core_052 = cgp_core_038 | input_g[1];
  assign cgp_core_054 = input_b[0] & input_a[0];
  assign cgp_core_057_not = ~input_f[1];
  assign cgp_core_058 = input_f[0] & input_c[1];
  assign cgp_core_060 = ~cgp_core_052;
  assign cgp_core_061 = input_a[0] & input_d[1];
  assign cgp_core_062 = cgp_core_051 ^ input_c[1];
  assign cgp_core_063 = ~(input_b[1] & input_f[1]);
  assign cgp_core_064 = ~(input_c[0] | input_a[0]);
  assign cgp_core_065 = ~(input_a[1] | input_g[1]);
  assign cgp_core_066 = ~(input_g[1] | cgp_core_063);
  assign cgp_core_068 = input_b[1] ^ cgp_core_063;
  assign cgp_core_069 = input_b[0] ^ input_f[1];
  assign cgp_core_070 = input_e[0] & input_b[0];
  assign cgp_core_071 = cgp_core_070 & input_d[1];
  assign cgp_core_072 = ~(input_f[0] & cgp_core_057_not);
  assign cgp_core_074 = input_d[1] | input_c[0];
  assign cgp_core_075 = input_d[1] & input_e[0];
  assign cgp_core_076 = input_e[0] & input_g[0];
  assign cgp_core_078 = input_e[0] & input_b[1];
  assign cgp_core_079 = input_f[0] | cgp_core_066;
  assign cgp_core_081 = input_b[1] | input_g[1];
  assign cgp_core_082 = input_e[1] | input_c[1];

  assign cgp_out[0] = 1'b1;
endmodule