module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;

  assign cgp_core_014 = input_f[0] & input_d[1];
  assign cgp_core_015 = input_c[1] ^ input_c[1];
  assign cgp_core_018 = input_d[1] & input_b[1];
  assign cgp_core_019 = ~(input_d[1] & input_a[0]);
  assign cgp_core_022 = ~(input_d[1] | input_a[1]);
  assign cgp_core_024 = ~input_f[1];
  assign cgp_core_025_not = ~input_d[0];
  assign cgp_core_026 = ~(input_a[0] | input_b[1]);
  assign cgp_core_031 = input_c[0] | input_c[0];
  assign cgp_core_034 = ~(input_e[1] | input_c[0]);
  assign cgp_core_035 = ~input_c[0];
  assign cgp_core_038 = ~input_b[0];
  assign cgp_core_039 = input_f[1] | input_a[1];
  assign cgp_core_040 = ~input_a[0];
  assign cgp_core_043 = input_a[0] | cgp_core_039;
  assign cgp_core_046 = input_d[1] | cgp_core_043;
  assign cgp_core_047 = ~(input_a[0] & input_e[0]);
  assign cgp_core_048 = input_f[1] ^ input_f[1];
  assign cgp_core_049 = input_c[1] & input_c[0];
  assign cgp_core_050 = input_e[1] & input_d[1];
  assign cgp_core_052 = ~(input_f[1] ^ input_c[1]);
  assign cgp_core_053 = ~(input_a[1] | input_a[0]);
  assign cgp_core_054 = ~(input_b[0] ^ input_d[1]);
  assign cgp_core_057 = input_d[0] | input_b[1];
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_062 = ~(input_d[1] ^ input_d[1]);
  assign cgp_core_063 = input_e[0] & input_e[1];
  assign cgp_core_064 = input_e[1] | input_f[0];
  assign cgp_core_067 = ~(input_d[0] | input_c[0]);
  assign cgp_core_068 = cgp_core_058 | cgp_core_046;
  assign cgp_core_069 = input_c[1] | cgp_core_068;
  assign cgp_core_070 = input_f[0] | input_f[1];
  assign cgp_core_072 = cgp_core_069 | input_e[1];

  assign cgp_out[0] = cgp_core_072;
endmodule