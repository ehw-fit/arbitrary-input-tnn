module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_013_not;
  wire cgp_core_015;
  wire cgp_core_016_not;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_033;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_054;

  assign cgp_core_012 = ~(input_e[0] & input_c[0]);
  assign cgp_core_013_not = ~input_a[1];
  assign cgp_core_015 = input_a[0] | input_e[1];
  assign cgp_core_016_not = ~input_b[1];
  assign cgp_core_018 = input_b[1] | input_b[0];
  assign cgp_core_019 = ~(input_b[0] & input_a[1]);
  assign cgp_core_020 = ~input_d[1];
  assign cgp_core_021 = input_c[1] | input_e[1];
  assign cgp_core_022 = input_c[1] & input_e[1];
  assign cgp_core_023 = cgp_core_021 | cgp_core_020;
  assign cgp_core_024 = cgp_core_021 & cgp_core_020;
  assign cgp_core_025 = cgp_core_022 | cgp_core_024;
  assign cgp_core_026 = ~(input_a[1] ^ input_c[0]);
  assign cgp_core_027 = ~input_a[1];
  assign cgp_core_029 = input_a[1] & cgp_core_023;
  assign cgp_core_033 = cgp_core_025 | cgp_core_029;
  assign cgp_core_037 = ~cgp_core_033;
  assign cgp_core_038 = cgp_core_018 & cgp_core_037;
  assign cgp_core_040 = ~(input_e[0] | cgp_core_033);
  assign cgp_core_042 = ~(input_e[0] ^ input_b[1]);
  assign cgp_core_043 = input_a[1] ^ input_e[0];
  assign cgp_core_045 = ~input_d[1];
  assign cgp_core_046 = ~(input_c[0] | input_e[1]);
  assign cgp_core_047 = ~(input_a[1] | input_c[0]);
  assign cgp_core_048 = input_b[0] ^ input_c[0];
  assign cgp_core_049 = input_a[0] & input_d[0];
  assign cgp_core_054 = cgp_core_040 | cgp_core_038;

  assign cgp_out[0] = cgp_core_054;
endmodule