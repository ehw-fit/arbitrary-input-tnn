module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032_not;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051_not;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_014 = input_c[1] & input_d[0];
  assign cgp_core_015 = ~input_d[0];
  assign cgp_core_017 = input_d[0] ^ input_b[2];
  assign cgp_core_018 = input_b[0] | input_a[2];
  assign cgp_core_020 = ~input_a[1];
  assign cgp_core_021 = input_a[2] | input_b[2];
  assign cgp_core_022 = input_a[2] & input_b[2];
  assign cgp_core_024 = input_a[1] & input_b[1];
  assign cgp_core_025 = cgp_core_022 | cgp_core_024;
  assign cgp_core_026 = ~input_b[2];
  assign cgp_core_028 = ~(input_b[2] & input_d[0]);
  assign cgp_core_029 = input_c[0] & input_c[2];
  assign cgp_core_030 = input_a[2] | input_b[2];
  assign cgp_core_032_not = ~input_a[2];
  assign cgp_core_036 = ~input_d[2];
  assign cgp_core_038 = ~input_d[2];
  assign cgp_core_039 = cgp_core_025 & cgp_core_038;
  assign cgp_core_040_not = ~input_a[2];
  assign cgp_core_041 = ~input_c[2];
  assign cgp_core_042 = cgp_core_021 & cgp_core_041;
  assign cgp_core_044 = input_a[0] & input_b[0];
  assign cgp_core_045 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_046 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_047 = ~(input_c[0] ^ input_c[1]);
  assign cgp_core_051_not = ~input_d[2];
  assign cgp_core_055 = input_a[1] ^ input_d[0];
  assign cgp_core_056 = input_d[1] ^ input_c[0];
  assign cgp_core_058 = cgp_core_042 | cgp_core_039;
  assign cgp_core_059 = ~input_c[1];

  assign cgp_out[0] = cgp_core_058;
endmodule