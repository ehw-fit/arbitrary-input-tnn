module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038_not;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_086;
  wire cgp_core_087_not;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_091_not;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_095;

  assign cgp_core_018 = ~(input_b[0] & input_f[1]);
  assign cgp_core_020 = ~(input_d[1] | input_b[0]);
  assign cgp_core_023 = ~(input_e[1] & input_e[1]);
  assign cgp_core_024 = input_a[1] | input_g[0];
  assign cgp_core_026 = input_a[0] & input_c[0];
  assign cgp_core_027 = ~(input_a[1] & input_e[1]);
  assign cgp_core_028 = input_a[1] & input_f[0];
  assign cgp_core_030 = input_f[1] & cgp_core_026;
  assign cgp_core_031 = cgp_core_028 | input_h[0];
  assign cgp_core_032 = ~input_a[0];
  assign cgp_core_033 = input_c[1] & input_d[0];
  assign cgp_core_035 = input_f[0] & input_e[0];
  assign cgp_core_036 = ~(input_b[0] & input_h[1]);
  assign cgp_core_038_not = ~input_g[1];
  assign cgp_core_039 = ~(cgp_core_036 ^ input_h[0]);
  assign cgp_core_042 = ~(input_g[0] | input_a[1]);
  assign cgp_core_044 = input_c[0] & cgp_core_038_not;
  assign cgp_core_045 = input_f[0] ^ cgp_core_042;
  assign cgp_core_046 = ~(input_h[1] | cgp_core_042);
  assign cgp_core_047 = input_c[1] & input_e[0];
  assign cgp_core_048 = input_b[1] | input_e[0];
  assign cgp_core_052 = input_a[1] ^ input_h[1];
  assign cgp_core_054 = input_c[0] | input_h[0];
  assign cgp_core_055 = ~(input_g[0] ^ input_f[0]);
  assign cgp_core_057 = input_d[0] | input_e[0];
  assign cgp_core_058 = input_g[0] ^ input_a[0];
  assign cgp_core_062 = ~(input_b[0] & input_h[1]);
  assign cgp_core_063 = ~(input_f[1] | input_a[1]);
  assign cgp_core_069 = ~(input_e[1] | input_f[1]);
  assign cgp_core_070 = ~(input_d[1] & input_f[1]);
  assign cgp_core_071 = cgp_core_069 & input_c[0];
  assign cgp_core_072 = input_d[0] & input_b[1];
  assign cgp_core_073 = ~input_a[1];
  assign cgp_core_076 = input_g[1] | input_b[1];
  assign cgp_core_077 = cgp_core_076 & input_g[1];
  assign cgp_core_078 = input_f[0] | input_a[1];
  assign cgp_core_079 = input_h[1] ^ cgp_core_078;
  assign cgp_core_080 = cgp_core_079 & input_c[0];
  assign cgp_core_082 = input_c[0] & input_h[1];
  assign cgp_core_083 = cgp_core_071 & input_h[1];
  assign cgp_core_084 = ~input_e[0];
  assign cgp_core_086 = ~(input_f[0] ^ input_h[1]);
  assign cgp_core_087_not = ~cgp_core_082;
  assign cgp_core_088 = ~(input_c[0] & input_a[1]);
  assign cgp_core_089 = ~(input_d[0] & cgp_core_088);
  assign cgp_core_091_not = ~input_b[1];
  assign cgp_core_092 = ~(input_f[1] & cgp_core_087_not);
  assign cgp_core_093 = ~(input_a[1] & input_b[0]);
  assign cgp_core_095 = input_c[0] | input_d[1];

  assign cgp_out[0] = 1'b1;
endmodule