module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_060_not;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_072;
  wire cgp_core_077_not;
  wire cgp_core_078;

  assign cgp_core_018 = input_a[0] & input_b[0];
  assign cgp_core_024 = ~input_d[1];
  assign cgp_core_026 = ~cgp_core_024;
  assign cgp_core_029 = input_d[2] ^ input_e[0];
  assign cgp_core_031 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_033 = input_a[0] | input_d[0];
  assign cgp_core_034 = input_e[2] ^ input_d[0];
  assign cgp_core_037 = ~(input_d[2] ^ input_a[1]);
  assign cgp_core_044 = input_e[2] & input_d[0];
  assign cgp_core_045 = ~(input_b[2] & input_b[2]);
  assign cgp_core_048 = input_c[2] | input_a[0];
  assign cgp_core_049 = input_c[2] & input_e[2];
  assign cgp_core_051 = ~(input_b[2] ^ input_c[2]);
  assign cgp_core_052 = input_b[1] | input_a[0];
  assign cgp_core_054 = input_b[1] & cgp_core_052;
  assign cgp_core_057 = ~(input_e[0] & input_c[1]);
  assign cgp_core_060_not = ~input_a[2];
  assign cgp_core_063 = ~(input_b[1] | input_c[2]);
  assign cgp_core_064 = cgp_core_063 | input_c[2];
  assign cgp_core_066 = ~(input_b[1] ^ input_d[1]);
  assign cgp_core_067 = ~cgp_core_045;
  assign cgp_core_069 = ~(input_e[1] | input_b[1]);
  assign cgp_core_072 = input_e[0] & input_c[0];
  assign cgp_core_077_not = ~input_a[1];
  assign cgp_core_078 = input_c[2] | input_d[0];

  assign cgp_out[0] = 1'b0;
endmodule