module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060_not;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_071;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_089;
  wire cgp_core_091;
  wire cgp_core_092_not;
  wire cgp_core_093;

  assign cgp_core_018 = ~input_d[0];
  assign cgp_core_021 = input_d[1] & input_h[1];
  assign cgp_core_023 = input_d[1] & input_c[1];
  assign cgp_core_026 = input_a[0] & input_e[0];
  assign cgp_core_027 = input_a[1] ^ input_d[0];
  assign cgp_core_028 = ~input_f[0];
  assign cgp_core_030 = ~(input_e[0] ^ cgp_core_026);
  assign cgp_core_032 = ~(input_a[0] | input_e[0]);
  assign cgp_core_034 = ~(input_b[0] ^ input_c[1]);
  assign cgp_core_035 = ~(input_a[0] & input_a[1]);
  assign cgp_core_037 = input_c[0] ^ input_c[1];
  assign cgp_core_039 = ~(input_f[0] | cgp_core_035);
  assign cgp_core_040 = cgp_core_037 | cgp_core_039;
  assign cgp_core_042 = input_f[0] | input_g[1];
  assign cgp_core_044 = input_f[1] & input_g[1];
  assign cgp_core_046 = input_e[0] & input_f[1];
  assign cgp_core_048 = ~(input_g[1] & input_a[1]);
  assign cgp_core_051 = ~input_e[1];
  assign cgp_core_057 = cgp_core_034 & cgp_core_048;
  assign cgp_core_059 = ~(input_h[0] | input_e[1]);
  assign cgp_core_060_not = ~input_a[0];
  assign cgp_core_061 = cgp_core_059 ^ input_a[0];
  assign cgp_core_062 = ~(input_e[1] & input_a[1]);
  assign cgp_core_063 = input_e[1] | cgp_core_062;
  assign cgp_core_066 = input_f[0] | input_h[0];
  assign cgp_core_067 = input_c[1] & cgp_core_063;
  assign cgp_core_071 = ~input_d[0];
  assign cgp_core_077 = input_h[1] & input_g[0];
  assign cgp_core_078 = ~cgp_core_066;
  assign cgp_core_080 = ~(input_f[1] & input_f[0]);
  assign cgp_core_083 = ~cgp_core_061;
  assign cgp_core_085 = ~input_e[0];
  assign cgp_core_086 = ~(input_a[1] | input_e[0]);
  assign cgp_core_089 = input_d[1] & input_h[0];
  assign cgp_core_091 = ~(input_b[0] ^ input_f[0]);
  assign cgp_core_092_not = ~cgp_core_091;
  assign cgp_core_093 = cgp_core_085 ^ cgp_core_080;

  assign cgp_out[0] = 1'b0;
endmodule