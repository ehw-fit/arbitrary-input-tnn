module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073_not;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_d[2] | input_a[0]);
  assign cgp_core_018 = ~input_b[1];
  assign cgp_core_019 = input_d[1] & input_b[1];
  assign cgp_core_022 = ~input_a[1];
  assign cgp_core_024 = ~(input_d[0] ^ input_b[1]);
  assign cgp_core_026 = ~input_a[1];
  assign cgp_core_028 = ~(input_c[0] & input_e[1]);
  assign cgp_core_030 = ~(input_d[0] & input_b[2]);
  assign cgp_core_031 = input_c[2] | input_a[0];
  assign cgp_core_032 = input_b[2] & input_a[2];
  assign cgp_core_034 = input_d[0] | input_d[0];
  assign cgp_core_035_not = ~input_b[2];
  assign cgp_core_036 = input_b[0] & input_c[1];
  assign cgp_core_037 = input_a[2] ^ input_e[1];
  assign cgp_core_038 = ~input_a[1];
  assign cgp_core_039 = ~(input_c[1] | input_b[0]);
  assign cgp_core_040 = input_c[2] | input_e[2];
  assign cgp_core_042 = input_b[2] & cgp_core_040;
  assign cgp_core_048 = ~(input_c[0] | input_a[0]);
  assign cgp_core_049 = input_d[1] | input_a[1];
  assign cgp_core_050 = input_a[2] | input_d[2];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_052 = ~(input_a[0] | input_a[2]);
  assign cgp_core_053 = cgp_core_050 & cgp_core_049;
  assign cgp_core_054 = cgp_core_051 | cgp_core_053;
  assign cgp_core_055 = input_d[1] | input_d[1];
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_064 = ~input_c[0];
  assign cgp_core_066 = input_c[2] | input_e[1];
  assign cgp_core_067 = input_c[2] ^ input_b[1];
  assign cgp_core_068 = input_d[2] & input_b[2];
  assign cgp_core_070 = ~(input_b[2] | input_b[1]);
  assign cgp_core_072 = ~input_d[1];
  assign cgp_core_073_not = ~input_d[0];
  assign cgp_core_074 = input_b[1] & input_d[1];
  assign cgp_core_075 = input_c[2] & input_e[2];
  assign cgp_core_076 = ~(input_d[0] | input_d[0]);
  assign cgp_core_077 = ~(input_d[2] ^ input_a[0]);
  assign cgp_core_078 = cgp_core_042 | cgp_core_075;
  assign cgp_core_079 = cgp_core_056 | cgp_core_078;

  assign cgp_out[0] = cgp_core_079;
endmodule