module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_010;
  wire cgp_core_011;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_043;

  assign cgp_core_010 = input_a[0] ^ input_a[1];
  assign cgp_core_011 = ~input_b[0];
  assign cgp_core_016 = ~(input_c[0] ^ input_d[0]);
  assign cgp_core_018 = ~(input_c[0] ^ input_c[1]);
  assign cgp_core_019 = input_b[1] | input_d[1];
  assign cgp_core_023 = ~(input_a[1] & input_c[1]);
  assign cgp_core_024_not = ~input_d[0];
  assign cgp_core_026 = input_d[0] | input_b[0];
  assign cgp_core_027 = input_b[0] | input_a[0];
  assign cgp_core_028 = ~(input_c[1] & input_d[1]);
  assign cgp_core_029 = ~input_c[1];
  assign cgp_core_030 = ~(input_a[0] | input_c[0]);
  assign cgp_core_033 = ~input_a[1];
  assign cgp_core_035 = ~(input_d[1] & input_a[0]);
  assign cgp_core_036 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_040 = cgp_core_033 | cgp_core_019;
  assign cgp_core_041 = ~input_b[1];
  assign cgp_core_042_not = ~input_d[1];
  assign cgp_core_043 = cgp_core_040 | input_c[1];

  assign cgp_out[0] = cgp_core_043;
endmodule