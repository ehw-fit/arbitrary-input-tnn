module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_014 = input_c[0] & input_b[0];
  assign cgp_core_015 = input_c[0] & input_f[0];
  assign cgp_core_017 = ~(input_e[0] ^ input_f[1]);
  assign cgp_core_018 = input_a[1] | cgp_core_015;
  assign cgp_core_019 = ~(input_c[0] | input_f[1]);
  assign cgp_core_020 = ~(input_f[1] ^ input_c[1]);
  assign cgp_core_021 = input_b[0] ^ input_f[0];
  assign cgp_core_025 = ~(input_b[0] & input_c[0]);
  assign cgp_core_027 = input_d[0] | input_c[1];
  assign cgp_core_028 = input_e[0] & input_b[1];
  assign cgp_core_029 = ~(input_d[1] | input_c[0]);
  assign cgp_core_031 = input_e[0] & input_d[1];
  assign cgp_core_033 = input_a[0] & input_d[0];
  assign cgp_core_034 = input_d[1] | cgp_core_033;
  assign cgp_core_035 = input_a[1] | cgp_core_034;
  assign cgp_core_036 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_037 = input_a[1] ^ input_d[0];
  assign cgp_core_038 = input_c[0] ^ input_d[1];
  assign cgp_core_040 = ~input_c[1];
  assign cgp_core_042 = ~(input_c[0] | input_b[0]);
  assign cgp_core_043 = ~(input_c[1] ^ input_b[1]);
  assign cgp_core_044 = input_c[1] | cgp_core_035;
  assign cgp_core_047 = ~input_b[0];
  assign cgp_core_048 = ~input_d[1];
  assign cgp_core_052 = ~(input_c[0] | input_d[1]);
  assign cgp_core_053 = input_c[1] & input_e[0];
  assign cgp_core_054 = ~(input_f[1] & input_d[1]);
  assign cgp_core_056 = ~(input_a[0] ^ input_d[1]);
  assign cgp_core_058 = ~input_d[0];
  assign cgp_core_061 = ~input_b[1];
  assign cgp_core_064_not = ~input_e[0];
  assign cgp_core_065 = ~(input_c[0] & input_c[1]);
  assign cgp_core_066 = ~(input_a[1] | input_c[1]);
  assign cgp_core_068 = cgp_core_018 | cgp_core_044;
  assign cgp_core_069 = input_e[1] | cgp_core_068;
  assign cgp_core_070 = input_c[1] | cgp_core_061;
  assign cgp_core_071 = input_f[1] | cgp_core_070;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;

  assign cgp_out[0] = cgp_core_072;
endmodule