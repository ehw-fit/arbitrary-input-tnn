module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063_not;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_095;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_101_not;
  wire cgp_core_103;
  wire cgp_core_106;
  wire cgp_core_110;

  assign cgp_core_020 = ~input_h[0];
  assign cgp_core_021 = input_e[0] ^ input_i[0];
  assign cgp_core_022 = ~(input_g[1] | input_g[0]);
  assign cgp_core_023 = input_h[1] & input_i[1];
  assign cgp_core_024 = ~(input_e[1] | input_i[1]);
  assign cgp_core_028 = ~input_b[0];
  assign cgp_core_030 = ~(input_e[1] & input_h[0]);
  assign cgp_core_032 = ~(input_e[0] | input_g[1]);
  assign cgp_core_033 = input_g[1] & input_f[0];
  assign cgp_core_034 = input_d[0] & input_d[1];
  assign cgp_core_036 = input_i[1] & input_g[1];
  assign cgp_core_038 = input_g[0] & input_b[1];
  assign cgp_core_039 = input_h[0] & input_b[0];
  assign cgp_core_042 = ~(input_g[0] & input_i[1]);
  assign cgp_core_044 = input_f[1] & input_a[1];
  assign cgp_core_046 = input_d[0] ^ input_a[0];
  assign cgp_core_047 = ~(input_a[0] ^ input_c[0]);
  assign cgp_core_048_not = ~input_d[0];
  assign cgp_core_049 = ~(input_f[1] & input_f[1]);
  assign cgp_core_050 = input_b[1] | input_a[1];
  assign cgp_core_054 = ~(input_a[0] ^ input_b[1]);
  assign cgp_core_055 = ~(input_c[0] & input_i[1]);
  assign cgp_core_056 = ~(input_g[1] | input_d[1]);
  assign cgp_core_058 = input_g[1] | input_f[1];
  assign cgp_core_059 = ~(input_f[0] ^ input_a[0]);
  assign cgp_core_060 = ~input_e[0];
  assign cgp_core_061 = input_e[1] & input_b[0];
  assign cgp_core_063_not = ~input_a[1];
  assign cgp_core_065 = input_e[1] | input_c[1];
  assign cgp_core_066 = cgp_core_058 | cgp_core_065;
  assign cgp_core_067 = cgp_core_058 & cgp_core_065;
  assign cgp_core_068 = ~(input_h[0] | input_e[1]);
  assign cgp_core_069 = ~(input_h[1] | input_e[1]);
  assign cgp_core_070 = input_e[1] | input_c[0];
  assign cgp_core_071 = ~(input_f[0] ^ input_a[1]);
  assign cgp_core_073 = input_b[0] & input_c[1];
  assign cgp_core_074 = ~input_g[1];
  assign cgp_core_075 = input_b[1] | cgp_core_066;
  assign cgp_core_076 = cgp_core_050 & cgp_core_066;
  assign cgp_core_078 = input_g[0] & input_c[0];
  assign cgp_core_079 = cgp_core_076 | cgp_core_078;
  assign cgp_core_081 = ~(input_f[1] ^ input_e[0]);
  assign cgp_core_082 = cgp_core_067 | cgp_core_079;
  assign cgp_core_084 = input_d[1] | input_b[1];
  assign cgp_core_085 = ~input_g[0];
  assign cgp_core_086 = ~(input_e[1] ^ input_d[0]);
  assign cgp_core_087 = ~cgp_core_082;
  assign cgp_core_088 = cgp_core_023 & cgp_core_087;
  assign cgp_core_091 = ~(input_c[1] & input_g[1]);
  assign cgp_core_092 = input_i[0] | input_a[1];
  assign cgp_core_093 = ~input_a[1];
  assign cgp_core_095 = ~(input_a[1] | cgp_core_075);
  assign cgp_core_097 = ~input_a[1];
  assign cgp_core_098 = ~input_e[0];
  assign cgp_core_099 = input_d[1] & cgp_core_095;
  assign cgp_core_100 = ~(input_c[0] | input_e[0]);
  assign cgp_core_101_not = ~input_e[0];
  assign cgp_core_103 = ~(input_f[1] & input_c[1]);
  assign cgp_core_106 = ~(input_a[0] | input_h[1]);
  assign cgp_core_110 = cgp_core_099 | cgp_core_088;

  assign cgp_out[0] = cgp_core_110;
endmodule