module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_054_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;

  assign cgp_core_014 = input_a[0] ^ input_b[1];
  assign cgp_core_015 = ~(input_b[1] ^ input_a[0]);
  assign cgp_core_018 = ~(input_d[0] ^ input_a[0]);
  assign cgp_core_019_not = ~input_d[0];
  assign cgp_core_021 = ~(input_d[1] & input_a[1]);
  assign cgp_core_022 = input_b[0] ^ input_e[0];
  assign cgp_core_023 = input_a[1] | input_e[1];
  assign cgp_core_025 = ~input_d[0];
  assign cgp_core_026 = ~(input_c[1] | cgp_core_022);
  assign cgp_core_027 = input_a[0] & input_b[1];
  assign cgp_core_028 = input_d[0] | input_f[0];
  assign cgp_core_029 = ~input_a[0];
  assign cgp_core_031 = ~(input_f[0] | input_d[1]);
  assign cgp_core_032 = ~(input_e[1] | input_c[0]);
  assign cgp_core_034 = ~(input_f[0] | input_c[1]);
  assign cgp_core_035 = ~cgp_core_027;
  assign cgp_core_036 = ~(input_d[0] & input_e[0]);
  assign cgp_core_039 = cgp_core_018 ^ cgp_core_032;
  assign cgp_core_042 = cgp_core_039 | input_d[0];
  assign cgp_core_044 = ~(input_a[1] | input_c[0]);
  assign cgp_core_045 = input_a[1] ^ input_d[0];
  assign cgp_core_046 = ~cgp_core_044;
  assign cgp_core_049 = cgp_core_036 | input_a[0];
  assign cgp_core_051 = input_b[1] ^ input_a[1];
  assign cgp_core_054_not = ~input_b[1];
  assign cgp_core_056 = input_a[1] | input_a[1];
  assign cgp_core_057 = input_a[1] ^ input_d[0];
  assign cgp_core_058 = ~input_c[0];
  assign cgp_core_059 = ~(input_c[1] ^ input_b[1]);
  assign cgp_core_060 = ~input_d[1];
  assign cgp_core_062 = input_f[1] & cgp_core_057;
  assign cgp_core_064 = cgp_core_028 & input_c[0];
  assign cgp_core_066 = ~input_f[1];
  assign cgp_core_067 = ~(cgp_core_066 | input_a[0]);
  assign cgp_core_069 = ~(input_a[1] | input_c[0]);
  assign cgp_core_070 = input_b[0] | input_b[1];
  assign cgp_core_071 = input_a[1] | input_a[0];

  assign cgp_out[0] = 1'b1;
endmodule