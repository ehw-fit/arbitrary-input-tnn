module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_065;

  assign cgp_core_017 = ~(input_d[0] | input_a[1]);
  assign cgp_core_018 = input_b[0] ^ input_c[0];
  assign cgp_core_020 = input_c[0] ^ input_d[0];
  assign cgp_core_021 = ~(input_f[0] & input_c[1]);
  assign cgp_core_022_not = ~input_a[0];
  assign cgp_core_023 = input_b[1] | input_d[1];
  assign cgp_core_024 = input_f[0] & input_d[1];
  assign cgp_core_025 = cgp_core_023 | input_e[1];
  assign cgp_core_026 = cgp_core_023 & input_d[0];
  assign cgp_core_027 = cgp_core_024 | cgp_core_026;
  assign cgp_core_028 = ~input_d[0];
  assign cgp_core_031 = input_e[1] & input_f[1];
  assign cgp_core_032 = input_b[0] | input_e[1];
  assign cgp_core_033 = input_b[1] & input_e[0];
  assign cgp_core_034 = cgp_core_031 | cgp_core_033;
  assign cgp_core_035 = input_c[1] | input_f[1];
  assign cgp_core_036 = input_f[0] ^ input_d[0];
  assign cgp_core_038 = cgp_core_025 & cgp_core_032;
  assign cgp_core_039 = ~(input_a[0] ^ input_f[1]);
  assign cgp_core_040 = ~(input_e[1] | input_a[1]);
  assign cgp_core_042 = cgp_core_027 | cgp_core_034;
  assign cgp_core_044 = input_f[1] | cgp_core_038;
  assign cgp_core_047 = ~(input_b[0] | input_c[0]);
  assign cgp_core_048 = ~cgp_core_042;
  assign cgp_core_049 = ~cgp_core_044;
  assign cgp_core_050 = input_a[1] & cgp_core_049;
  assign cgp_core_051 = cgp_core_050 & cgp_core_048;
  assign cgp_core_052 = ~(input_a[1] ^ cgp_core_044);
  assign cgp_core_053 = cgp_core_052 & cgp_core_048;
  assign cgp_core_057 = ~(input_b[1] & input_c[0]);
  assign cgp_core_058 = input_c[1] & cgp_core_053;
  assign cgp_core_059 = input_e[1] ^ input_d[1];
  assign cgp_core_061 = ~input_b[1];
  assign cgp_core_062 = input_b[0] & input_e[0];
  assign cgp_core_063 = input_c[1] & cgp_core_058;
  assign cgp_core_064_not = ~input_f[0];
  assign cgp_core_065 = cgp_core_051 | cgp_core_063;

  assign cgp_out[0] = cgp_core_065;
endmodule