module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_038_not;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_074;

  assign cgp_core_017 = input_b[0] ^ input_c[0];
  assign cgp_core_018 = input_b[0] & input_c[0];
  assign cgp_core_019 = ~(input_b[1] & input_d[1]);
  assign cgp_core_020 = input_b[1] & input_c[1];
  assign cgp_core_021 = cgp_core_019 ^ cgp_core_018;
  assign cgp_core_022 = cgp_core_019 & cgp_core_018;
  assign cgp_core_023 = cgp_core_020 | cgp_core_022;
  assign cgp_core_025 = ~input_b[2];
  assign cgp_core_027 = input_b[2] & cgp_core_023;
  assign cgp_core_028 = input_c[2] | cgp_core_027;
  assign cgp_core_029 = input_d[0] ^ input_c[2];
  assign cgp_core_030 = input_d[0] & input_e[0];
  assign cgp_core_031 = input_d[1] & input_e[1];
  assign cgp_core_032 = input_d[1] & input_b[1];
  assign cgp_core_033 = cgp_core_031 ^ cgp_core_030;
  assign cgp_core_034 = input_d[2] & cgp_core_030;
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038_not = ~input_c[1];
  assign cgp_core_042 = input_d[1] & input_a[2];
  assign cgp_core_043 = cgp_core_021 ^ cgp_core_033;
  assign cgp_core_044 = cgp_core_021 & cgp_core_033;
  assign cgp_core_045 = ~cgp_core_043;
  assign cgp_core_046 = ~(cgp_core_043 | input_a[0]);
  assign cgp_core_047 = cgp_core_044 | cgp_core_046;
  assign cgp_core_050_not = ~cgp_core_047;
  assign cgp_core_051 = input_e[2] & cgp_core_047;
  assign cgp_core_052 = input_d[1] | cgp_core_051;
  assign cgp_core_055 = input_b[2] ^ cgp_core_052;
  assign cgp_core_056 = input_b[0] & input_c[1];
  assign cgp_core_057 = input_b[2] | input_d[0];
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = ~input_e[1];
  assign cgp_core_060 = ~cgp_core_055;
  assign cgp_core_061 = ~input_e[1];
  assign cgp_core_062 = cgp_core_061 & cgp_core_059;
  assign cgp_core_063 = ~input_d[0];
  assign cgp_core_064 = input_a[2] & input_a[0];
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066 = ~(input_a[2] ^ cgp_core_050_not);
  assign cgp_core_068 = ~input_b[0];
  assign cgp_core_069 = input_a[2] & cgp_core_068;
  assign cgp_core_071 = ~(input_a[1] ^ cgp_core_045);
  assign cgp_core_074 = input_a[0] & input_c[0];

  assign cgp_out[0] = 1'b0;
endmodule