module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052_not;
  wire cgp_core_053;

  assign cgp_core_013 = input_b[1] | input_c[1];
  assign cgp_core_014 = input_c[0] & input_c[0];
  assign cgp_core_016 = input_b[0] & input_e[1];
  assign cgp_core_017 = ~(input_a[0] | input_e[1]);
  assign cgp_core_020 = input_a[0] & input_c[1];
  assign cgp_core_022 = ~(input_b[0] & cgp_core_016);
  assign cgp_core_023 = ~(input_a[0] ^ input_b[1]);
  assign cgp_core_024 = input_a[0] | input_b[0];
  assign cgp_core_025 = cgp_core_022 & input_e[0];
  assign cgp_core_026 = input_a[0] ^ cgp_core_025;
  assign cgp_core_029 = input_c[1] & input_a[0];
  assign cgp_core_032 = ~input_b[0];
  assign cgp_core_035_not = ~input_a[0];
  assign cgp_core_036 = input_c[0] & input_d[0];
  assign cgp_core_037 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_039 = ~(input_d[1] ^ input_a[1]);
  assign cgp_core_040 = ~(input_a[1] & input_c[1]);
  assign cgp_core_042 = ~(input_c[0] | input_c[1]);
  assign cgp_core_043 = ~cgp_core_042;
  assign cgp_core_045 = ~(input_d[1] | input_c[1]);
  assign cgp_core_046 = ~input_b[1];
  assign cgp_core_047 = input_b[1] & input_a[0];
  assign cgp_core_048 = input_c[0] | cgp_core_045;
  assign cgp_core_051 = ~(input_a[1] ^ input_e[1]);
  assign cgp_core_052_not = ~input_b[1];
  assign cgp_core_053 = input_a[0] | input_c[0];

  assign cgp_out[0] = input_a[1];
endmodule