module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_030;
  wire cgp_core_031_not;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_014 = ~(input_b[2] ^ input_d[2]);
  assign cgp_core_016 = ~(input_d[1] & input_c[2]);
  assign cgp_core_018 = ~input_b[0];
  assign cgp_core_019 = ~input_d[1];
  assign cgp_core_020 = ~(input_b[1] | input_b[1]);
  assign cgp_core_021 = ~input_a[2];
  assign cgp_core_025 = input_d[2] | input_d[0];
  assign cgp_core_028 = ~input_b[0];
  assign cgp_core_029_not = ~input_a[0];
  assign cgp_core_030 = ~(input_c[1] & input_a[2]);
  assign cgp_core_031_not = ~input_b[0];
  assign cgp_core_034 = ~(input_b[1] ^ input_d[0]);
  assign cgp_core_037 = ~(input_c[0] | input_c[0]);
  assign cgp_core_038 = ~input_d[2];
  assign cgp_core_039 = input_a[2] & cgp_core_038;
  assign cgp_core_040 = input_a[0] ^ input_a[2];
  assign cgp_core_041_not = ~input_c[1];
  assign cgp_core_042 = ~(input_d[0] & input_d[0]);
  assign cgp_core_044 = ~(input_c[1] & input_a[0]);
  assign cgp_core_045 = input_a[0] ^ input_d[2];
  assign cgp_core_049 = ~input_a[2];
  assign cgp_core_051 = input_d[2] | input_c[1];
  assign cgp_core_052 = input_c[2] ^ input_d[2];
  assign cgp_core_053 = input_a[1] ^ input_c[2];
  assign cgp_core_055 = ~(input_c[2] ^ input_c[2]);
  assign cgp_core_056 = ~(input_c[1] ^ input_d[2]);
  assign cgp_core_058 = input_b[2] | cgp_core_039;
  assign cgp_core_059 = ~(input_a[1] | input_b[2]);

  assign cgp_out[0] = cgp_core_058;
endmodule