module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018_not;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_082;

  assign cgp_core_016 = input_e[1] | input_c[0];
  assign cgp_core_017 = ~(input_a[0] | input_c[0]);
  assign cgp_core_018_not = ~input_a[0];
  assign cgp_core_020 = ~(input_d[0] & input_f[0]);
  assign cgp_core_021 = ~input_e[0];
  assign cgp_core_022 = ~(input_a[0] | input_a[1]);
  assign cgp_core_023 = input_e[0] | input_g[0];
  assign cgp_core_024 = input_e[0] & input_g[0];
  assign cgp_core_025 = input_e[1] | input_b[0];
  assign cgp_core_026 = ~(input_f[1] & input_g[1]);
  assign cgp_core_028 = input_d[1] & cgp_core_024;
  assign cgp_core_029 = cgp_core_026 | cgp_core_028;
  assign cgp_core_031 = input_b[1] & cgp_core_023;
  assign cgp_core_032 = ~(input_d[1] & input_c[1]);
  assign cgp_core_035 = cgp_core_032 & cgp_core_031;
  assign cgp_core_038 = input_d[1] & input_g[0];
  assign cgp_core_039 = cgp_core_016 ^ input_a[1];
  assign cgp_core_042 = cgp_core_020 & input_b[0];
  assign cgp_core_046 = input_e[0] | input_c[1];
  assign cgp_core_048 = cgp_core_046 ^ input_b[1];
  assign cgp_core_049 = ~cgp_core_046;
  assign cgp_core_051 = cgp_core_038 ^ cgp_core_049;
  assign cgp_core_052 = cgp_core_038 & cgp_core_049;
  assign cgp_core_053_not = ~input_b[0];
  assign cgp_core_054 = input_b[0] & input_f[0];
  assign cgp_core_055 = input_b[0] ^ input_f[1];
  assign cgp_core_056 = ~input_g[0];
  assign cgp_core_057 = cgp_core_055 & cgp_core_054;
  assign cgp_core_058 = input_f[0] & cgp_core_054;
  assign cgp_core_059 = input_c[0] & input_c[1];
  assign cgp_core_060 = ~(cgp_core_052 | cgp_core_052);
  assign cgp_core_061 = cgp_core_051 | cgp_core_060;
  assign cgp_core_062 = ~cgp_core_051;
  assign cgp_core_063 = ~(cgp_core_062 | input_c[0]);
  assign cgp_core_064 = ~input_e[1];
  assign cgp_core_065 = cgp_core_048 & cgp_core_064;
  assign cgp_core_068 = cgp_core_048 & input_c[1];
  assign cgp_core_069 = ~cgp_core_057;
  assign cgp_core_070 = ~(input_d[0] ^ cgp_core_069);
  assign cgp_core_072 = ~(input_d[0] ^ cgp_core_057);
  assign cgp_core_076 = input_f[0] & input_d[0];
  assign cgp_core_077 = ~cgp_core_039;
  assign cgp_core_082 = input_e[0] | input_b[1];

  assign cgp_out[0] = 1'b1;
endmodule