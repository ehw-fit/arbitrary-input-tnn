module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_039_not;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = input_a[0] ^ input_e[0];
  assign cgp_core_018 = input_b[0] ^ input_d[1];
  assign cgp_core_019 = input_c[1] ^ input_e[0];
  assign cgp_core_020 = ~(input_e[1] & cgp_core_017);
  assign cgp_core_021 = cgp_core_018 ^ input_c[1];
  assign cgp_core_024 = ~(input_b[0] & input_g[0]);
  assign cgp_core_026 = input_e[1] | input_g[1];
  assign cgp_core_027_not = ~cgp_core_024;
  assign cgp_core_028_not = ~cgp_core_024;
  assign cgp_core_029 = input_d[0] ^ cgp_core_028_not;
  assign cgp_core_039_not = ~input_f[1];
  assign cgp_core_041_not = ~input_g[1];
  assign cgp_core_042 = input_b[0] ^ input_f[0];
  assign cgp_core_043 = input_b[0] & input_e[0];
  assign cgp_core_046 = ~(input_a[1] | input_g[0]);
  assign cgp_core_047 = input_c[1] & input_f[0];
  assign cgp_core_049_not = ~cgp_core_042;
  assign cgp_core_050 = input_a[0] & input_g[0];
  assign cgp_core_051 = ~(input_d[0] | input_g[1]);
  assign cgp_core_052 = input_d[0] & input_c[0];
  assign cgp_core_053 = ~(input_b[1] & cgp_core_050);
  assign cgp_core_054 = cgp_core_051 & cgp_core_050;
  assign cgp_core_055 = cgp_core_052 & input_b[0];
  assign cgp_core_058 = ~input_a[1];
  assign cgp_core_059 = ~(cgp_core_041_not & cgp_core_058);
  assign cgp_core_060 = ~(input_d[0] & input_c[1]);
  assign cgp_core_061 = ~input_d[1];
  assign cgp_core_063 = input_c[0] & input_g[1];
  assign cgp_core_064_not = ~input_f[1];
  assign cgp_core_066 = ~input_g[0];
  assign cgp_core_068 = input_a[1] & input_c[0];
  assign cgp_core_069 = ~(input_a[1] ^ input_c[1]);
  assign cgp_core_070 = input_c[1] & input_a[0];
  assign cgp_core_071 = cgp_core_049_not ^ cgp_core_049_not;
  assign cgp_core_072 = input_d[0] & cgp_core_071;
  assign cgp_core_073 = cgp_core_072 | input_f[0];
  assign cgp_core_074 = input_g[1] | input_a[1];
  assign cgp_core_075 = cgp_core_074 & cgp_core_070;
  assign cgp_core_077 = cgp_core_059 | input_f[0];
  assign cgp_core_078 = ~(cgp_core_063 & input_b[0]);
  assign cgp_core_079 = input_e[0] | input_c[1];

  assign cgp_out[0] = 1'b1;
endmodule