module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_021_not;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_035;
  wire cgp_core_039_not;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051_not;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_b[0] | input_d[2]);
  assign cgp_core_020 = ~(input_c[1] & input_c[1]);
  assign cgp_core_021_not = ~input_a[0];
  assign cgp_core_023 = input_e[2] ^ input_c[1];
  assign cgp_core_025 = ~(input_b[2] ^ input_a[0]);
  assign cgp_core_026 = input_e[2] ^ input_a[1];
  assign cgp_core_027 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_028 = ~(input_d[0] & input_b[2]);
  assign cgp_core_029_not = ~input_c[2];
  assign cgp_core_030 = ~(input_d[1] | input_d[2]);
  assign cgp_core_033 = input_d[1] & input_d[1];
  assign cgp_core_034_not = ~input_c[1];
  assign cgp_core_035 = input_d[1] ^ input_e[1];
  assign cgp_core_039_not = ~input_a[1];
  assign cgp_core_042 = ~(input_e[0] | input_c[0]);
  assign cgp_core_043_not = ~input_b[2];
  assign cgp_core_044 = input_c[2] | input_d[2];
  assign cgp_core_048 = ~(input_d[1] | input_a[0]);
  assign cgp_core_049 = ~(input_b[2] & input_d[1]);
  assign cgp_core_050 = ~(input_c[1] | input_e[0]);
  assign cgp_core_051_not = ~input_c[1];
  assign cgp_core_052 = ~input_b[0];
  assign cgp_core_053 = ~input_e[0];
  assign cgp_core_054 = input_e[0] ^ input_c[2];
  assign cgp_core_056 = ~(input_d[1] & input_a[2]);
  assign cgp_core_057 = input_b[0] | input_b[1];
  assign cgp_core_058 = input_a[1] & input_a[0];
  assign cgp_core_060 = input_e[2] ^ input_a[1];
  assign cgp_core_061 = ~(input_b[2] ^ input_d[0]);
  assign cgp_core_063 = ~(input_d[2] ^ input_a[2]);
  assign cgp_core_065 = input_b[1] ^ input_c[1];
  assign cgp_core_067 = ~(input_d[0] ^ input_a[1]);
  assign cgp_core_068 = input_d[1] & input_a[0];
  assign cgp_core_070 = ~(input_c[2] ^ input_a[0]);
  assign cgp_core_072 = input_b[1] | input_e[0];
  assign cgp_core_073 = input_a[0] | input_e[0];
  assign cgp_core_074 = ~(input_c[2] & input_a[1]);
  assign cgp_core_075 = ~(input_d[1] | input_c[2]);
  assign cgp_core_077 = input_e[1] | input_d[2];
  assign cgp_core_079 = ~(input_a[2] ^ input_e[1]);

  assign cgp_out[0] = 1'b0;
endmodule