module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_014_not;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_027_not;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047_not;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;

  assign cgp_core_012 = input_d[1] | input_d[0];
  assign cgp_core_014_not = ~input_c[0];
  assign cgp_core_019 = input_b[1] ^ input_a[0];
  assign cgp_core_021 = input_a[1] & input_b[0];
  assign cgp_core_022 = ~input_b[1];
  assign cgp_core_027_not = ~input_c[1];
  assign cgp_core_029 = ~(input_e[0] ^ input_d[1]);
  assign cgp_core_030 = ~(input_d[0] ^ input_a[0]);
  assign cgp_core_031 = input_e[1] | input_d[1];
  assign cgp_core_033 = input_e[1] | input_c[1];
  assign cgp_core_034 = ~(input_a[1] ^ input_b[0]);
  assign cgp_core_035 = ~(input_e[0] | input_b[0]);
  assign cgp_core_037 = ~cgp_core_033;
  assign cgp_core_038 = input_b[1] & cgp_core_037;
  assign cgp_core_040 = ~(input_a[1] | input_a[0]);
  assign cgp_core_042 = ~(input_c[0] ^ input_c[1]);
  assign cgp_core_043 = ~(input_c[0] & input_c[1]);
  assign cgp_core_046 = input_b[0] & cgp_core_040;
  assign cgp_core_047_not = ~input_d[0];
  assign cgp_core_048 = ~(input_c[0] ^ input_d[1]);
  assign cgp_core_049 = ~(input_d[0] ^ input_c[1]);
  assign cgp_core_051 = input_d[1] & cgp_core_046;
  assign cgp_core_052 = input_b[1] | input_a[1];
  assign cgp_core_053 = cgp_core_038 | cgp_core_051;

  assign cgp_out[0] = cgp_core_053;
endmodule