module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049_not;
  wire cgp_core_051;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_066;

  assign cgp_core_014 = ~(input_a[1] & input_b[1]);
  assign cgp_core_015 = ~(input_e[1] & input_f[1]);
  assign cgp_core_017 = input_a[1] & input_c[1];
  assign cgp_core_018 = ~(input_e[1] ^ input_a[1]);
  assign cgp_core_022 = ~(input_a[1] | input_e[1]);
  assign cgp_core_023 = input_c[1] ^ input_d[1];
  assign cgp_core_024 = ~(input_a[1] & input_c[0]);
  assign cgp_core_025 = ~(input_f[1] ^ input_c[0]);
  assign cgp_core_026 = input_e[1] ^ input_c[0];
  assign cgp_core_030 = ~(input_b[1] | input_f[0]);
  assign cgp_core_033 = ~(input_e[1] & input_b[1]);
  assign cgp_core_034 = ~(input_e[0] & input_b[1]);
  assign cgp_core_035 = input_b[0] & input_a[0];
  assign cgp_core_036 = ~(input_b[0] ^ input_b[1]);
  assign cgp_core_037 = input_a[0] ^ input_a[1];
  assign cgp_core_038 = ~(input_e[0] & input_c[0]);
  assign cgp_core_040 = input_e[1] | input_e[0];
  assign cgp_core_041 = input_e[0] ^ input_f[0];
  assign cgp_core_042 = ~(input_e[1] | input_c[1]);
  assign cgp_core_045 = input_c[0] ^ input_c[0];
  assign cgp_core_046 = input_d[1] | input_b[1];
  assign cgp_core_047 = ~input_d[1];
  assign cgp_core_048 = ~cgp_core_046;
  assign cgp_core_049_not = ~input_b[1];
  assign cgp_core_051 = cgp_core_017 & cgp_core_048;
  assign cgp_core_055 = input_c[0] & input_b[0];
  assign cgp_core_056 = ~(input_a[0] | input_f[1]);
  assign cgp_core_057 = input_a[1] ^ input_f[1];
  assign cgp_core_058 = ~(input_a[0] | input_e[1]);
  assign cgp_core_059 = ~(input_d[0] & input_c[1]);
  assign cgp_core_060 = ~(input_f[1] & input_c[1]);
  assign cgp_core_064 = input_d[0] ^ input_d[1];
  assign cgp_core_066 = ~(input_d[0] & input_b[0]);

  assign cgp_out[0] = cgp_core_051;
endmodule