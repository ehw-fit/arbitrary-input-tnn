module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042_not;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_053;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062_not;

  assign cgp_core_015 = input_a[0] & input_c[0];
  assign cgp_core_016 = input_f[1] ^ input_c[1];
  assign cgp_core_017 = input_a[1] & input_c[1];
  assign cgp_core_018 = input_d[0] ^ cgp_core_015;
  assign cgp_core_021 = ~input_b[0];
  assign cgp_core_024 = ~input_a[1];
  assign cgp_core_025 = input_d[1] ^ input_d[0];
  assign cgp_core_028 = input_e[0] & input_f[0];
  assign cgp_core_030 = input_f[0] ^ input_e[1];
  assign cgp_core_035 = cgp_core_021 ^ input_b[1];
  assign cgp_core_037 = cgp_core_025 ^ input_f[1];
  assign cgp_core_038 = cgp_core_025 & input_f[0];
  assign cgp_core_039 = ~(input_a[1] | input_e[0]);
  assign cgp_core_040 = input_f[0] & input_b[0];
  assign cgp_core_042_not = ~input_f[1];
  assign cgp_core_047 = ~input_f[1];
  assign cgp_core_048 = ~input_a[0];
  assign cgp_core_053 = cgp_core_017 & input_f[1];
  assign cgp_core_057 = cgp_core_018 ^ cgp_core_039;
  assign cgp_core_059 = ~input_e[1];
  assign cgp_core_060 = input_d[1] | cgp_core_059;
  assign cgp_core_062_not = ~cgp_core_035;

  assign cgp_out[0] = 1'b0;
endmodule