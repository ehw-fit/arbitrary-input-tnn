module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_050;
  wire cgp_core_054_not;
  wire cgp_core_059;

  assign cgp_core_015 = input_b[2] | input_c[2];
  assign cgp_core_016_not = ~input_d[1];
  assign cgp_core_017 = input_d[1] & input_b[2];
  assign cgp_core_018 = input_a[1] | input_a[0];
  assign cgp_core_019_not = ~input_c[1];
  assign cgp_core_021 = ~(input_b[2] | input_a[1]);
  assign cgp_core_024 = ~(input_a[2] ^ input_a[1]);
  assign cgp_core_025 = input_b[0] | input_d[0];
  assign cgp_core_026 = ~input_c[2];
  assign cgp_core_027 = input_a[2] ^ input_a[2];
  assign cgp_core_028 = ~input_b[2];
  assign cgp_core_030 = ~input_c[0];
  assign cgp_core_032 = input_c[2] ^ input_c[1];
  assign cgp_core_034 = input_c[0] | input_b[1];
  assign cgp_core_036 = ~(input_c[0] ^ input_a[1]);
  assign cgp_core_037 = input_c[1] | input_d[2];
  assign cgp_core_038 = input_b[0] | input_d[0];
  assign cgp_core_040 = ~input_c[2];
  assign cgp_core_041 = input_c[0] & input_c[1];
  assign cgp_core_043 = input_a[2] & cgp_core_040;
  assign cgp_core_044 = input_b[1] & input_d[0];
  assign cgp_core_045 = ~(input_c[0] | input_d[1]);
  assign cgp_core_050 = ~(input_c[0] ^ input_b[2]);
  assign cgp_core_054_not = ~input_d[2];
  assign cgp_core_059 = input_b[2] | cgp_core_043;

  assign cgp_out[0] = cgp_core_059;
endmodule