module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_017;
  wire cgp_core_019_not;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033_not;
  wire cgp_core_036_not;
  wire cgp_core_037;
  wire cgp_core_038_not;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;

  assign cgp_core_011 = ~(input_c[1] ^ input_a[0]);
  assign cgp_core_012 = ~(input_c[1] ^ input_a[0]);
  assign cgp_core_017 = input_c[1] & input_a[0];
  assign cgp_core_019_not = ~input_d[1];
  assign cgp_core_021 = ~(input_a[1] ^ input_c[0]);
  assign cgp_core_024 = input_a[1] ^ input_a[0];
  assign cgp_core_025 = ~input_a[1];
  assign cgp_core_029 = input_d[1] ^ input_a[1];
  assign cgp_core_030 = ~input_a[1];
  assign cgp_core_033_not = ~input_c[0];
  assign cgp_core_036_not = ~input_d[1];
  assign cgp_core_037 = ~(input_b[0] | input_d[0]);
  assign cgp_core_038_not = ~input_a[1];
  assign cgp_core_039 = ~(input_c[1] | input_a[0]);
  assign cgp_core_040 = input_c[1] | cgp_core_030;
  assign cgp_core_042 = input_d[1] | input_b[1];
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;

  assign cgp_out[0] = cgp_core_043;
endmodule