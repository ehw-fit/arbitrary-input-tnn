module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_078;

  assign cgp_core_017 = input_b[0] ^ input_b[2];
  assign cgp_core_018 = input_b[1] & input_a[2];
  assign cgp_core_019 = input_b[1] ^ input_c[1];
  assign cgp_core_020 = input_d[1] & input_c[1];
  assign cgp_core_022 = cgp_core_019 & cgp_core_018;
  assign cgp_core_023 = ~(input_e[0] & cgp_core_022);
  assign cgp_core_024 = input_b[2] ^ input_c[2];
  assign cgp_core_025 = input_c[1] & input_c[2];
  assign cgp_core_027 = input_e[0] ^ cgp_core_023;
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_029 = input_a[1] ^ input_e[0];
  assign cgp_core_031 = input_d[1] ^ input_e[1];
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_035 = cgp_core_032 | input_c[1];
  assign cgp_core_036 = input_d[2] ^ input_e[2];
  assign cgp_core_037 = ~(input_d[2] & input_d[2]);
  assign cgp_core_038 = cgp_core_036 ^ cgp_core_035;
  assign cgp_core_041 = ~(cgp_core_017 & input_a[0]);
  assign cgp_core_042 = ~(cgp_core_017 ^ input_b[0]);
  assign cgp_core_043 = cgp_core_019 & cgp_core_031;
  assign cgp_core_044 = cgp_core_019 & input_b[0];
  assign cgp_core_046 = cgp_core_043 & cgp_core_042;
  assign cgp_core_047 = ~(cgp_core_044 ^ cgp_core_046);
  assign cgp_core_050 = input_a[0] ^ cgp_core_047;
  assign cgp_core_051 = ~(input_e[2] | cgp_core_047);
  assign cgp_core_052 = ~input_e[2];
  assign cgp_core_054 = cgp_core_028 & input_c[1];
  assign cgp_core_057 = input_b[0] | input_a[1];
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = ~input_b[1];
  assign cgp_core_060 = ~cgp_core_052;
  assign cgp_core_061 = ~input_e[2];
  assign cgp_core_062 = input_e[0] & cgp_core_059;
  assign cgp_core_063 = input_c[2] | cgp_core_050;
  assign cgp_core_064 = input_b[0] & input_b[1];
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066 = input_b[2] & cgp_core_050;
  assign cgp_core_071 = ~(input_a[1] ^ input_a[0]);
  assign cgp_core_073 = ~cgp_core_041;
  assign cgp_core_076 = ~(input_a[0] & input_e[2]);
  assign cgp_core_078 = ~(input_c[2] ^ cgp_core_065);

  assign cgp_out[0] = 1'b0;
endmodule