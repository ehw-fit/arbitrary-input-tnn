module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028_not;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040_not;
  wire cgp_core_041;
  wire cgp_core_042;

  assign cgp_core_012 = input_a[0] | input_a[0];
  assign cgp_core_013 = ~input_a[0];
  assign cgp_core_014 = ~input_c[2];
  assign cgp_core_017 = ~(input_c[0] ^ input_b[1]);
  assign cgp_core_019 = input_c[0] ^ input_b[0];
  assign cgp_core_022 = ~input_c[1];
  assign cgp_core_023 = ~input_c[1];
  assign cgp_core_025 = ~input_a[2];
  assign cgp_core_026 = ~(input_c[2] | input_a[2]);
  assign cgp_core_028_not = ~input_a[1];
  assign cgp_core_030 = input_b[2] | input_b[2];
  assign cgp_core_033 = ~(input_b[0] & input_c[1]);
  assign cgp_core_035 = input_c[2] ^ input_a[0];
  assign cgp_core_038 = ~input_c[1];
  assign cgp_core_039 = input_c[2] ^ input_a[0];
  assign cgp_core_040_not = ~input_a[0];
  assign cgp_core_041 = ~input_a[0];
  assign cgp_core_042 = ~(input_a[1] ^ input_c[2]);

  assign cgp_out[0] = cgp_core_026;
endmodule