module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052_not;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_089;
  wire cgp_core_096;

  assign cgp_core_018 = input_d[0] | input_h[0];
  assign cgp_core_019 = input_d[0] & input_h[0];
  assign cgp_core_020 = ~input_h[1];
  assign cgp_core_021 = input_d[1] & input_h[1];
  assign cgp_core_023 = input_a[0] | input_b[0];
  assign cgp_core_026 = input_a[0] & cgp_core_018;
  assign cgp_core_027 = input_b[0] | input_c[1];
  assign cgp_core_028 = input_a[1] & cgp_core_019;
  assign cgp_core_029 = ~(input_a[0] & input_d[1]);
  assign cgp_core_030 = input_a[1] & cgp_core_026;
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = cgp_core_021 | cgp_core_031;
  assign cgp_core_033 = cgp_core_021 & cgp_core_031;
  assign cgp_core_043 = ~(input_h[1] ^ input_b[1]);
  assign cgp_core_045 = ~(input_b[0] & input_d[0]);
  assign cgp_core_046 = input_h[1] ^ input_h[0];
  assign cgp_core_047 = input_f[0] | input_f[1];
  assign cgp_core_049 = ~(input_b[1] | input_g[1]);
  assign cgp_core_050 = input_h[1] & input_f[1];
  assign cgp_core_051 = ~(input_b[0] | input_f[1]);
  assign cgp_core_052_not = ~input_h[0];
  assign cgp_core_054_not = ~input_b[0];
  assign cgp_core_055 = input_f[0] ^ input_f[1];
  assign cgp_core_056 = input_h[1] & input_f[1];
  assign cgp_core_057 = input_c[0] | input_e[0];
  assign cgp_core_060 = input_c[0] | input_g[1];
  assign cgp_core_061 = input_b[0] & input_d[1];
  assign cgp_core_063 = ~(input_a[1] | input_c[1]);
  assign cgp_core_066 = ~(input_h[1] ^ input_a[0]);
  assign cgp_core_067 = ~(input_b[0] & input_a[1]);
  assign cgp_core_068 = input_f[1] | input_g[0];
  assign cgp_core_069 = input_e[1] | input_f[1];
  assign cgp_core_071 = input_e[1] ^ input_h[0];
  assign cgp_core_072 = ~input_g[1];
  assign cgp_core_073 = input_a[0] | input_d[0];
  assign cgp_core_075 = cgp_core_033 & cgp_core_072;
  assign cgp_core_076 = ~(input_b[1] | cgp_core_069);
  assign cgp_core_080 = cgp_core_032 & cgp_core_076;
  assign cgp_core_082 = input_d[0] ^ input_g[1];
  assign cgp_core_084 = ~(input_g[0] & input_h[1]);
  assign cgp_core_085 = ~(input_h[1] | input_g[1]);
  assign cgp_core_089 = ~(input_g[0] & input_h[0]);
  assign cgp_core_096 = cgp_core_080 | cgp_core_075;

  assign cgp_out[0] = cgp_core_096;
endmodule