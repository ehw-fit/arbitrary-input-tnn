module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;

  assign cgp_core_020 = input_f[2] ^ input_b[0];
  assign cgp_core_021 = input_a[0] & input_b[0];
  assign cgp_core_022 = input_a[1] ^ input_b[1];
  assign cgp_core_023 = input_a[2] & input_b[1];
  assign cgp_core_024 = cgp_core_022 ^ input_c[1];
  assign cgp_core_025 = cgp_core_022 & input_b[0];
  assign cgp_core_026 = cgp_core_023 | cgp_core_025;
  assign cgp_core_027 = input_f[2] ^ input_f[2];
  assign cgp_core_028 = input_a[2] & input_b[2];
  assign cgp_core_029 = ~input_a[1];
  assign cgp_core_030 = input_c[1] & cgp_core_026;
  assign cgp_core_033 = input_c[0] & input_f[0];
  assign cgp_core_034 = input_b[2] ^ input_d[1];
  assign cgp_core_035 = input_c[1] & input_d[1];
  assign cgp_core_036 = ~(cgp_core_034 | input_f[2]);
  assign cgp_core_037 = cgp_core_034 & cgp_core_033;
  assign cgp_core_038 = input_f[0] | cgp_core_037;
  assign cgp_core_039 = input_c[2] & input_d[2];
  assign cgp_core_040 = input_c[2] & input_d[2];
  assign cgp_core_041 = cgp_core_039 ^ cgp_core_038;
  assign cgp_core_042 = cgp_core_039 & cgp_core_038;
  assign cgp_core_043 = cgp_core_040 | input_d[1];
  assign cgp_core_044 = input_e[0] | input_e[1];
  assign cgp_core_045 = input_e[0] & input_f[0];
  assign cgp_core_046 = input_e[1] ^ input_f[1];
  assign cgp_core_047 = input_e[1] & input_f[1];
  assign cgp_core_049 = input_d[0] & cgp_core_045;
  assign cgp_core_050 = cgp_core_047 | cgp_core_049;
  assign cgp_core_051 = input_e[2] ^ input_f[2];
  assign cgp_core_052 = input_e[2] & input_f[2];
  assign cgp_core_053 = cgp_core_051 ^ input_d[1];
  assign cgp_core_054 = input_c[1] & input_b[0];
  assign cgp_core_055 = ~cgp_core_052;
  assign cgp_core_056 = ~(input_d[1] | cgp_core_044);
  assign cgp_core_058 = cgp_core_036 ^ input_f[1];
  assign cgp_core_059 = cgp_core_036 & cgp_core_046;
  assign cgp_core_060 = cgp_core_058 ^ cgp_core_044;
  assign cgp_core_061 = cgp_core_058 & cgp_core_044;
  assign cgp_core_062 = cgp_core_059 | cgp_core_061;
  assign cgp_core_063 = cgp_core_041 ^ cgp_core_053;
  assign cgp_core_064 = cgp_core_041 & cgp_core_053;
  assign cgp_core_065 = ~(cgp_core_063 ^ input_d[2]);
  assign cgp_core_066 = cgp_core_063 & cgp_core_062;
  assign cgp_core_067 = input_c[1] | input_c[0];
  assign cgp_core_068 = cgp_core_043 ^ cgp_core_055;
  assign cgp_core_069 = cgp_core_043 & cgp_core_055;
  assign cgp_core_070 = cgp_core_068 ^ cgp_core_067;
  assign cgp_core_071 = cgp_core_068 & input_a[1];
  assign cgp_core_072 = ~(cgp_core_069 & cgp_core_071);
  assign cgp_core_073 = ~cgp_core_072;
  assign cgp_core_074 = ~cgp_core_072;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = input_f[1] & cgp_core_075;
  assign cgp_core_077 = cgp_core_076 & input_e[2];
  assign cgp_core_078 = ~(input_f[1] ^ cgp_core_070);
  assign cgp_core_079 = input_e[2] & cgp_core_074;
  assign cgp_core_080 = ~input_a[2];
  assign cgp_core_081 = ~(cgp_core_029 | input_f[0]);
  assign cgp_core_085 = ~cgp_core_060;
  assign cgp_core_086 = cgp_core_024 & cgp_core_085;
  assign cgp_core_090 = ~input_b[1];
  assign cgp_core_091 = cgp_core_020 & input_c[2];
  assign cgp_core_093 = ~(cgp_core_020 ^ cgp_core_056);

  assign cgp_out[0] = 1'b0;
endmodule