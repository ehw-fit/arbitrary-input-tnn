module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023_not;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061_not;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_072;

  assign cgp_core_014 = input_e[1] ^ input_f[1];
  assign cgp_core_017 = ~(input_a[1] | input_b[1]);
  assign cgp_core_018 = ~input_b[0];
  assign cgp_core_019 = input_d[0] & input_f[0];
  assign cgp_core_020 = input_c[1] | cgp_core_019;
  assign cgp_core_021 = ~(input_f[1] | input_e[0]);
  assign cgp_core_022 = ~(input_e[0] | input_d[0]);
  assign cgp_core_023_not = ~input_b[0];
  assign cgp_core_025 = ~(input_d[1] | input_b[0]);
  assign cgp_core_027 = input_b[1] & input_b[0];
  assign cgp_core_028 = ~(input_c[1] | input_d[1]);
  assign cgp_core_029 = ~(input_d[1] | input_c[0]);
  assign cgp_core_030 = ~(input_e[0] | input_c[1]);
  assign cgp_core_035 = input_f[1] | input_d[1];
  assign cgp_core_036 = ~(input_d[1] ^ input_e[0]);
  assign cgp_core_037 = ~(input_c[0] & input_a[1]);
  assign cgp_core_042 = input_a[0] & input_c[0];
  assign cgp_core_043 = input_e[1] | cgp_core_042;
  assign cgp_core_044 = cgp_core_020 | cgp_core_035;
  assign cgp_core_046 = cgp_core_044 | cgp_core_043;
  assign cgp_core_048 = ~(input_b[0] | input_c[0]);
  assign cgp_core_054 = ~(input_e[1] ^ input_f[1]);
  assign cgp_core_056 = ~(input_e[0] ^ input_d[1]);
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_061_not = ~input_c[0];
  assign cgp_core_064 = input_c[0] ^ input_d[0];
  assign cgp_core_065 = input_f[1] ^ input_d[0];
  assign cgp_core_068 = cgp_core_058 | cgp_core_046;
  assign cgp_core_069 = input_a[1] | cgp_core_068;
  assign cgp_core_072 = input_d[1] & input_d[0];

  assign cgp_out[0] = cgp_core_069;
endmodule