module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_034;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[0] | input_a[2];
  assign cgp_core_016_not = ~input_a[10];
  assign cgp_core_017 = ~(input_a[5] & input_a[11]);
  assign cgp_core_018 = input_a[9] | input_a[6];
  assign cgp_core_022 = input_a[6] & input_a[5];
  assign cgp_core_025_not = ~input_a[0];
  assign cgp_core_026 = input_a[3] ^ input_a[4];
  assign cgp_core_027 = ~(input_a[1] & input_a[5]);
  assign cgp_core_028 = ~(input_a[5] ^ input_a[5]);
  assign cgp_core_030 = input_a[11] ^ input_a[4];
  assign cgp_core_034 = ~(input_a[0] | input_a[3]);
  assign cgp_core_038 = ~(input_a[10] & input_a[4]);
  assign cgp_core_039 = input_a[3] & input_a[7];
  assign cgp_core_041 = ~input_a[11];
  assign cgp_core_042 = input_a[3] ^ input_a[6];
  assign cgp_core_043_not = ~input_a[3];
  assign cgp_core_044 = ~(input_a[5] | input_a[11]);
  assign cgp_core_045 = input_a[3] & input_a[7];
  assign cgp_core_051 = ~(input_a[6] ^ input_a[3]);
  assign cgp_core_053 = ~input_a[10];
  assign cgp_core_064 = ~input_a[0];
  assign cgp_core_065 = ~input_a[0];
  assign cgp_core_066 = ~(input_a[11] & input_a[5]);
  assign cgp_core_067 = ~input_a[2];
  assign cgp_core_070 = input_a[2] | input_a[4];
  assign cgp_core_073 = input_a[5] ^ input_a[4];
  assign cgp_core_074 = input_a[1] & input_a[9];
  assign cgp_core_075 = ~(input_a[1] ^ input_a[9]);
  assign cgp_core_076 = input_a[2] ^ input_a[5];
  assign cgp_core_077 = input_a[5] & input_a[5];
  assign cgp_core_078 = input_a[1] & input_a[8];

  assign cgp_out[0] = input_a[3];
  assign cgp_out[1] = 1'b0;
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = input_a[6];
endmodule