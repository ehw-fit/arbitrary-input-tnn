module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_063;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_080_not;

  assign cgp_core_017 = input_e[1] | input_d[1];
  assign cgp_core_018 = input_c[1] ^ input_c[0];
  assign cgp_core_020 = ~(input_e[2] ^ input_c[2]);
  assign cgp_core_023 = ~(input_c[0] | input_b[0]);
  assign cgp_core_025 = ~(input_b[2] & input_a[2]);
  assign cgp_core_027 = ~(input_d[2] & input_a[2]);
  assign cgp_core_028 = input_b[2] | input_a[2];
  assign cgp_core_029_not = ~input_c[0];
  assign cgp_core_032 = input_d[1] & input_c[1];
  assign cgp_core_033 = input_a[1] | input_e[0];
  assign cgp_core_034 = ~(input_b[1] | input_b[0]);
  assign cgp_core_036 = input_d[2] | input_e[2];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038 = cgp_core_036 | cgp_core_032;
  assign cgp_core_039 = cgp_core_036 & cgp_core_032;
  assign cgp_core_040 = cgp_core_037 | cgp_core_039;
  assign cgp_core_043 = input_c[2] & input_d[2];
  assign cgp_core_045 = input_e[0] | input_d[0];
  assign cgp_core_046 = ~(input_b[2] | input_b[0]);
  assign cgp_core_048 = input_d[2] ^ input_a[2];
  assign cgp_core_049 = input_c[2] & cgp_core_038;
  assign cgp_core_050 = input_a[0] ^ input_a[2];
  assign cgp_core_053 = cgp_core_040 | cgp_core_049;
  assign cgp_core_056 = ~(input_c[1] ^ input_e[1]);
  assign cgp_core_057 = ~cgp_core_053;
  assign cgp_core_058 = cgp_core_028 & cgp_core_057;
  assign cgp_core_059 = input_e[0] ^ input_a[0];
  assign cgp_core_063 = input_e[0] & input_d[1];
  assign cgp_core_067 = input_a[1] ^ input_a[2];
  assign cgp_core_068 = input_b[1] ^ input_b[1];
  assign cgp_core_069 = input_e[2] ^ input_b[1];
  assign cgp_core_070 = ~(input_e[2] & input_e[1]);
  assign cgp_core_071 = input_e[2] ^ input_c[1];
  assign cgp_core_072 = input_e[0] ^ input_e[2];
  assign cgp_core_075 = ~input_d[1];
  assign cgp_core_076 = ~(input_e[0] & input_b[2]);
  assign cgp_core_080_not = ~input_c[0];

  assign cgp_out[0] = cgp_core_058;
endmodule