module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_069;
  wire cgp_core_071_not;
  wire cgp_core_076;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017 = input_e[2] & input_b[2];
  assign cgp_core_018 = input_a[2] ^ input_d[1];
  assign cgp_core_019 = ~(input_e[2] ^ input_c[2]);
  assign cgp_core_020 = ~(input_d[0] & input_c[0]);
  assign cgp_core_024 = input_a[0] & input_d[1];
  assign cgp_core_032 = ~(input_d[1] | input_c[2]);
  assign cgp_core_033 = ~(input_b[0] & input_d[2]);
  assign cgp_core_035 = input_d[0] & input_c[1];
  assign cgp_core_036 = ~(input_e[2] | input_c[2]);
  assign cgp_core_037 = ~input_d[1];
  assign cgp_core_038 = ~(input_e[1] ^ input_d[0]);
  assign cgp_core_041 = input_b[1] & input_a[2];
  assign cgp_core_045 = input_e[1] & input_b[2];
  assign cgp_core_048 = input_c[0] & input_b[0];
  assign cgp_core_049 = input_d[0] | input_e[2];
  assign cgp_core_050 = ~input_a[0];
  assign cgp_core_052 = ~(input_d[1] ^ input_e[0]);
  assign cgp_core_053 = ~(input_b[1] | input_a[0]);
  assign cgp_core_054 = ~(input_e[0] ^ input_e[0]);
  assign cgp_core_056 = input_b[0] ^ input_d[2];
  assign cgp_core_058 = ~input_d[2];
  assign cgp_core_060 = ~(input_c[1] & input_b[0]);
  assign cgp_core_061 = ~(input_a[0] & input_c[0]);
  assign cgp_core_062 = input_a[1] | input_a[0];
  assign cgp_core_063 = ~(input_a[0] | input_e[0]);
  assign cgp_core_064 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_069 = input_a[2] | input_a[1];
  assign cgp_core_071_not = ~input_a[0];
  assign cgp_core_076 = ~(input_e[2] ^ input_e[0]);
  assign cgp_core_079 = ~(input_c[0] | input_e[1]);
  assign cgp_core_080 = ~(input_d[1] ^ input_b[1]);

  assign cgp_out[0] = cgp_core_036;
endmodule