module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_082;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_097_not;
  wire cgp_core_099;
  wire cgp_core_101;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_110;

  assign cgp_core_020 = input_h[1] ^ input_f[1];
  assign cgp_core_021 = ~(input_h[0] ^ input_b[1]);
  assign cgp_core_022_not = ~input_f[1];
  assign cgp_core_023 = ~(input_h[1] ^ input_a[0]);
  assign cgp_core_024 = input_d[0] | input_a[1];
  assign cgp_core_025 = input_d[1] & input_g[1];
  assign cgp_core_027 = ~input_a[0];
  assign cgp_core_032 = ~(input_d[1] ^ input_b[0]);
  assign cgp_core_035 = ~input_f[1];
  assign cgp_core_036 = ~input_a[1];
  assign cgp_core_039 = ~input_i[1];
  assign cgp_core_041 = ~input_d[1];
  assign cgp_core_042 = input_c[1] | input_b[1];
  assign cgp_core_045 = ~(input_c[1] & input_d[1]);
  assign cgp_core_046 = input_c[0] | input_g[0];
  assign cgp_core_047 = input_c[1] ^ input_a[1];
  assign cgp_core_049 = input_a[1] | input_g[1];
  assign cgp_core_050 = cgp_core_042 | cgp_core_049;
  assign cgp_core_051 = cgp_core_042 & cgp_core_049;
  assign cgp_core_052 = input_a[0] ^ input_h[0];
  assign cgp_core_054_not = ~input_i[0];
  assign cgp_core_056 = ~(input_f[0] | input_i[0]);
  assign cgp_core_057 = input_c[0] & input_g[0];
  assign cgp_core_058 = input_e[1] | cgp_core_057;
  assign cgp_core_060 = input_i[0] | input_d[0];
  assign cgp_core_061 = input_g[1] ^ input_c[0];
  assign cgp_core_063 = input_h[0] | input_e[0];
  assign cgp_core_064 = input_h[0] | input_g[1];
  assign cgp_core_065 = ~(input_h[1] & input_c[1]);
  assign cgp_core_067 = ~(input_c[0] & input_a[1]);
  assign cgp_core_069 = ~(input_f[0] ^ input_d[1]);
  assign cgp_core_070 = ~(input_e[0] ^ input_d[0]);
  assign cgp_core_071 = ~(input_g[0] | input_d[0]);
  assign cgp_core_072 = ~(input_e[0] ^ input_h[0]);
  assign cgp_core_073 = ~input_c[0];
  assign cgp_core_075 = cgp_core_050 | cgp_core_058;
  assign cgp_core_076 = cgp_core_050 & cgp_core_058;
  assign cgp_core_078 = input_f[1] | input_e[1];
  assign cgp_core_082 = cgp_core_051 | cgp_core_076;
  assign cgp_core_086 = ~(input_i[1] & input_f[1]);
  assign cgp_core_087 = ~(input_g[1] | input_d[1]);
  assign cgp_core_089 = input_i[1] & input_c[0];
  assign cgp_core_090 = ~(input_f[1] | cgp_core_082);
  assign cgp_core_091 = cgp_core_090 & input_i[1];
  assign cgp_core_092 = ~(input_i[1] & input_i[0]);
  assign cgp_core_094 = input_h[1] & cgp_core_091;
  assign cgp_core_095 = ~(input_c[1] | cgp_core_075);
  assign cgp_core_097_not = ~input_f[0];
  assign cgp_core_099 = ~(input_e[1] & input_h[1]);
  assign cgp_core_101 = input_d[1] & cgp_core_095;
  assign cgp_core_104 = ~(input_g[1] & input_d[1]);
  assign cgp_core_105 = ~input_c[0];
  assign cgp_core_110 = cgp_core_094 | cgp_core_101;

  assign cgp_out[0] = cgp_core_110;
endmodule