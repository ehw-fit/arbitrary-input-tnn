module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032_not;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090_not;
  wire cgp_core_094;
  wire cgp_core_096;
  wire cgp_core_097_not;
  wire cgp_core_099;
  wire cgp_core_101;
  wire cgp_core_102;
  wire cgp_core_103;
  wire cgp_core_105;
  wire cgp_core_107;
  wire cgp_core_109;
  wire cgp_core_110;

  assign cgp_core_020 = ~(input_d[0] & input_h[1]);
  assign cgp_core_021 = input_b[0] & input_e[1];
  assign cgp_core_022 = input_h[1] | input_i[1];
  assign cgp_core_023 = input_h[1] & input_i[1];
  assign cgp_core_025 = input_b[1] ^ input_a[0];
  assign cgp_core_028 = ~(input_e[0] ^ input_f[1]);
  assign cgp_core_029 = input_a[1] & input_c[0];
  assign cgp_core_030 = input_d[1] & cgp_core_022;
  assign cgp_core_032_not = ~input_e[0];
  assign cgp_core_034 = cgp_core_023 | cgp_core_030;
  assign cgp_core_035 = ~input_a[1];
  assign cgp_core_036 = ~(input_h[1] | input_a[0]);
  assign cgp_core_037 = input_f[0] & input_b[0];
  assign cgp_core_038 = input_b[1] | input_c[1];
  assign cgp_core_039 = input_b[1] & input_c[1];
  assign cgp_core_040 = cgp_core_038 | cgp_core_037;
  assign cgp_core_041 = cgp_core_038 & cgp_core_037;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_043_not = ~input_i[1];
  assign cgp_core_044 = input_h[1] | input_a[0];
  assign cgp_core_045 = ~(input_c[1] | input_c[1]);
  assign cgp_core_046 = input_a[1] & cgp_core_040;
  assign cgp_core_047 = ~input_i[1];
  assign cgp_core_048 = ~(input_a[0] ^ input_g[0]);
  assign cgp_core_051 = input_a[1] & cgp_core_046;
  assign cgp_core_053 = input_g[1] | input_g[0];
  assign cgp_core_054 = ~(input_a[1] ^ input_c[0]);
  assign cgp_core_055 = ~input_h[0];
  assign cgp_core_057 = input_g[1] & input_h[1];
  assign cgp_core_058 = ~input_a[0];
  assign cgp_core_059 = input_b[0] ^ input_b[0];
  assign cgp_core_060 = input_b[1] & input_i[1];
  assign cgp_core_061 = input_e[1] | input_f[1];
  assign cgp_core_062 = input_e[1] & input_f[1];
  assign cgp_core_063 = ~input_c[1];
  assign cgp_core_064 = cgp_core_061 & input_g[1];
  assign cgp_core_065 = cgp_core_062 | cgp_core_064;
  assign cgp_core_066 = input_e[0] | input_i[0];
  assign cgp_core_068 = ~(input_e[1] & input_d[1]);
  assign cgp_core_069 = ~(input_h[1] | input_d[0]);
  assign cgp_core_070 = input_e[0] | input_h[0];
  assign cgp_core_071 = ~(input_e[1] ^ input_f[1]);
  assign cgp_core_072 = ~input_g[0];
  assign cgp_core_073 = ~(input_d[0] ^ input_i[1]);
  assign cgp_core_074 = ~(input_a[1] | input_d[1]);
  assign cgp_core_075 = input_d[1] & input_i[1];
  assign cgp_core_078 = input_d[0] | input_g[0];
  assign cgp_core_080 = cgp_core_051 | cgp_core_065;
  assign cgp_core_081 = ~(input_e[0] & input_i[0]);
  assign cgp_core_082 = cgp_core_080 | cgp_core_042;
  assign cgp_core_084 = input_f[0] ^ input_b[0];
  assign cgp_core_085 = input_c[0] ^ input_h[0];
  assign cgp_core_087 = input_d[0] | input_b[0];
  assign cgp_core_089 = ~(input_g[0] & input_h[0]);
  assign cgp_core_090_not = ~cgp_core_082;
  assign cgp_core_094 = input_c[1] ^ input_h[0];
  assign cgp_core_096 = cgp_core_034 & cgp_core_090_not;
  assign cgp_core_097_not = ~input_h[0];
  assign cgp_core_099 = ~(input_c[1] & input_h[1]);
  assign cgp_core_101 = ~(input_g[1] & input_a[0]);
  assign cgp_core_102 = input_g[0] ^ input_h[1];
  assign cgp_core_103 = ~(input_d[0] & input_f[1]);
  assign cgp_core_105 = ~(input_i[1] & input_f[0]);
  assign cgp_core_107 = ~input_h[0];
  assign cgp_core_109 = input_g[0] ^ input_a[0];
  assign cgp_core_110 = ~(input_b[1] | input_h[1]);

  assign cgp_out[0] = cgp_core_096;
endmodule