module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041_not;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;

  assign cgp_core_014 = ~(input_b[0] & input_a[1]);
  assign cgp_core_017 = ~input_e[1];
  assign cgp_core_018 = ~(input_b[0] & input_c[0]);
  assign cgp_core_020 = input_a[1] & input_c[1];
  assign cgp_core_023 = ~(input_c[0] | input_a[0]);
  assign cgp_core_025 = ~(input_b[0] | input_c[0]);
  assign cgp_core_028 = ~(input_b[1] & input_b[0]);
  assign cgp_core_030 = ~(input_b[1] | input_d[0]);
  assign cgp_core_031 = ~(input_f[0] & input_c[0]);
  assign cgp_core_032_not = ~input_c[0];
  assign cgp_core_033 = input_c[1] ^ input_d[0];
  assign cgp_core_038 = ~(input_d[1] ^ input_e[0]);
  assign cgp_core_039 = ~(input_b[1] | input_e[1]);
  assign cgp_core_041_not = ~input_a[1];
  assign cgp_core_045 = ~(input_f[0] & input_d[0]);
  assign cgp_core_046 = ~input_b[1];
  assign cgp_core_047 = input_f[1] ^ input_b[1];
  assign cgp_core_048 = ~input_d[1];
  assign cgp_core_050 = ~input_f[1];
  assign cgp_core_052 = input_d[0] ^ input_c[0];
  assign cgp_core_053 = input_c[1] & cgp_core_048;
  assign cgp_core_054 = ~input_f[1];
  assign cgp_core_055 = input_a[1] & cgp_core_054;
  assign cgp_core_056 = cgp_core_055 & cgp_core_053;
  assign cgp_core_057 = ~(input_c[0] ^ input_b[1]);
  assign cgp_core_058 = ~input_d[1];
  assign cgp_core_060 = input_c[0] & input_f[0];
  assign cgp_core_061 = input_f[0] ^ input_f[0];
  assign cgp_core_063 = ~(input_c[1] ^ input_c[0]);

  assign cgp_out[0] = cgp_core_056;
endmodule