module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020_not;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045_not;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_095;
  wire cgp_core_098;

  assign cgp_core_020_not = ~input_a[0];
  assign cgp_core_021 = ~(input_b[0] & input_b[0]);
  assign cgp_core_023 = input_b[1] | input_a[0];
  assign cgp_core_024 = ~(input_a[2] ^ input_f[1]);
  assign cgp_core_027 = input_a[2] ^ input_b[2];
  assign cgp_core_028 = ~(input_f[0] | input_a[0]);
  assign cgp_core_029 = ~input_f[0];
  assign cgp_core_031 = input_f[1] & input_d[1];
  assign cgp_core_032 = input_a[0] & input_d[0];
  assign cgp_core_033_not = ~input_d[0];
  assign cgp_core_034 = input_c[1] | input_a[0];
  assign cgp_core_036 = input_b[0] | input_b[2];
  assign cgp_core_037 = ~(cgp_core_034 ^ cgp_core_033_not);
  assign cgp_core_039 = ~(input_e[0] & input_d[2]);
  assign cgp_core_041 = ~(input_b[1] & input_f[0]);
  assign cgp_core_043 = input_e[2] | input_b[1];
  assign cgp_core_045_not = ~input_f[0];
  assign cgp_core_047 = input_c[0] | input_f[1];
  assign cgp_core_048 = input_d[0] ^ input_b[2];
  assign cgp_core_049 = ~input_b[1];
  assign cgp_core_051 = ~input_a[2];
  assign cgp_core_052 = input_c[2] ^ input_f[1];
  assign cgp_core_053 = cgp_core_051 & input_e[0];
  assign cgp_core_054 = ~(input_a[2] & input_c[1]);
  assign cgp_core_055 = input_d[1] | input_d[2];
  assign cgp_core_056 = input_f[0] ^ input_c[2];
  assign cgp_core_058 = ~(input_d[1] | input_b[2]);
  assign cgp_core_059 = cgp_core_036 & cgp_core_048;
  assign cgp_core_062 = ~input_d[2];
  assign cgp_core_063 = input_f[1] ^ input_d[0];
  assign cgp_core_064 = ~(input_b[0] | input_d[1]);
  assign cgp_core_065 = ~(input_c[2] & input_c[1]);
  assign cgp_core_066 = ~(input_a[2] & input_e[2]);
  assign cgp_core_068_not = ~input_b[2];
  assign cgp_core_070 = input_c[2] ^ input_c[0];
  assign cgp_core_071 = ~input_a[2];
  assign cgp_core_074 = ~input_f[2];
  assign cgp_core_075 = ~(input_a[1] & input_b[1]);
  assign cgp_core_077 = input_b[1] & input_f[1];
  assign cgp_core_078 = input_c[2] | input_a[0];
  assign cgp_core_079 = input_b[2] & input_a[2];
  assign cgp_core_080 = ~(input_e[0] ^ cgp_core_065);
  assign cgp_core_081 = ~input_e[2];
  assign cgp_core_082 = cgp_core_081 | input_f[1];
  assign cgp_core_086 = input_e[0] & input_e[1];
  assign cgp_core_088 = ~(input_b[2] | input_e[2]);
  assign cgp_core_092 = input_e[0] | input_b[0];
  assign cgp_core_093 = ~(input_f[0] ^ input_e[0]);
  assign cgp_core_095 = ~(input_a[2] & input_d[1]);
  assign cgp_core_098 = input_f[0] | input_b[0];

  assign cgp_out[0] = 1'b0;
endmodule