module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061_not;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_075_not;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079_not;
  wire cgp_core_080;
  wire cgp_core_081_not;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_091;
  wire cgp_core_093;

  assign cgp_core_018 = input_a[1] & input_e[1];
  assign cgp_core_019 = ~(input_d[1] ^ input_c[0]);
  assign cgp_core_022 = ~(input_a[0] | input_c[1]);
  assign cgp_core_023 = ~(input_h[0] & input_a[1]);
  assign cgp_core_024 = input_f[1] & input_f[0];
  assign cgp_core_026 = ~(input_g[0] & input_f[0]);
  assign cgp_core_027 = input_d[0] & cgp_core_022;
  assign cgp_core_029 = ~(input_b[1] | input_a[1]);
  assign cgp_core_031 = input_d[0] | input_f[1];
  assign cgp_core_033 = input_f[1] | input_b[0];
  assign cgp_core_034 = input_b[1] & input_d[1];
  assign cgp_core_036 = ~input_c[0];
  assign cgp_core_040 = input_a[0] & input_a[0];
  assign cgp_core_042 = ~(input_f[0] ^ input_b[1]);
  assign cgp_core_044 = ~(input_b[1] | input_c[0]);
  assign cgp_core_045_not = ~input_a[1];
  assign cgp_core_046 = ~input_f[0];
  assign cgp_core_048 = ~input_e[1];
  assign cgp_core_054 = input_c[0] | input_d[1];
  assign cgp_core_055 = input_a[0] & input_a[0];
  assign cgp_core_056 = input_f[1] & input_c[1];
  assign cgp_core_058 = input_e[1] | input_b[0];
  assign cgp_core_061_not = ~input_e[0];
  assign cgp_core_062 = ~(input_a[1] & cgp_core_058);
  assign cgp_core_063 = input_f[0] | input_a[0];
  assign cgp_core_065 = input_a[0] ^ input_a[0];
  assign cgp_core_067 = input_d[1] & input_h[0];
  assign cgp_core_068 = ~(input_h[1] ^ input_c[0]);
  assign cgp_core_070 = input_d[0] | input_e[0];
  assign cgp_core_071 = input_f[1] & input_d[1];
  assign cgp_core_075_not = ~input_h[1];
  assign cgp_core_076 = ~input_f[1];
  assign cgp_core_077 = input_b[1] | input_c[0];
  assign cgp_core_078 = input_a[1] | input_f[0];
  assign cgp_core_079_not = ~input_a[0];
  assign cgp_core_080 = ~(input_f[1] | input_a[0]);
  assign cgp_core_081_not = ~input_d[1];
  assign cgp_core_086 = ~(input_a[1] ^ input_d[1]);
  assign cgp_core_087 = ~input_b[1];
  assign cgp_core_089 = input_b[0] ^ input_b[0];
  assign cgp_core_091 = ~(input_h[0] | input_d[0]);
  assign cgp_core_093 = ~(input_b[1] | input_h[0]);

  assign cgp_out[0] = input_d[0];
endmodule