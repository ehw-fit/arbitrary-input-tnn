module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052_not;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_101;
  wire cgp_core_102;
  wire cgp_core_104;
  wire cgp_core_105_not;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_108;
  wire cgp_core_109;
  wire cgp_core_110;

  assign cgp_core_020 = input_h[0] ^ input_i[0];
  assign cgp_core_021 = input_h[0] & input_i[0];
  assign cgp_core_022 = input_h[1] ^ input_i[1];
  assign cgp_core_023 = input_h[1] & input_i[1];
  assign cgp_core_024 = cgp_core_022 ^ cgp_core_021;
  assign cgp_core_025 = cgp_core_022 & cgp_core_021;
  assign cgp_core_026 = cgp_core_023 | cgp_core_025;
  assign cgp_core_027 = input_d[0] ^ cgp_core_020;
  assign cgp_core_028 = input_d[0] & cgp_core_020;
  assign cgp_core_029 = input_d[1] ^ cgp_core_024;
  assign cgp_core_030 = input_d[1] & cgp_core_024;
  assign cgp_core_031 = cgp_core_029 ^ cgp_core_028;
  assign cgp_core_032 = cgp_core_029 & cgp_core_028;
  assign cgp_core_033 = cgp_core_030 | cgp_core_032;
  assign cgp_core_034 = cgp_core_026 ^ cgp_core_033;
  assign cgp_core_035 = cgp_core_026 & cgp_core_033;
  assign cgp_core_036 = input_b[0] ^ input_c[0];
  assign cgp_core_037 = input_b[0] & input_c[0];
  assign cgp_core_038 = input_b[1] ^ input_c[1];
  assign cgp_core_039 = input_b[1] & input_c[1];
  assign cgp_core_040 = cgp_core_038 ^ cgp_core_037;
  assign cgp_core_041 = cgp_core_038 & cgp_core_037;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_043 = input_a[0] ^ cgp_core_036;
  assign cgp_core_044 = input_a[0] & cgp_core_036;
  assign cgp_core_045 = input_a[1] ^ cgp_core_040;
  assign cgp_core_046 = input_a[1] & cgp_core_040;
  assign cgp_core_047 = cgp_core_045 ^ cgp_core_044;
  assign cgp_core_048 = cgp_core_045 & cgp_core_044;
  assign cgp_core_049 = cgp_core_046 | cgp_core_048;
  assign cgp_core_050 = cgp_core_042 | cgp_core_049;
  assign cgp_core_051 = cgp_core_042 & cgp_core_049;
  assign cgp_core_052_not = ~input_i[0];
  assign cgp_core_053 = input_f[0] & input_g[0];
  assign cgp_core_054 = input_f[1] ^ input_g[1];
  assign cgp_core_055 = input_f[1] & input_g[1];
  assign cgp_core_056 = cgp_core_054 ^ cgp_core_053;
  assign cgp_core_057 = cgp_core_054 & cgp_core_053;
  assign cgp_core_058 = cgp_core_055 | cgp_core_057;
  assign cgp_core_059 = ~input_e[0];
  assign cgp_core_060 = input_e[1] | input_h[1];
  assign cgp_core_061 = input_e[1] ^ cgp_core_056;
  assign cgp_core_062 = input_e[1] & cgp_core_056;
  assign cgp_core_063 = cgp_core_061 ^ input_e[0];
  assign cgp_core_064 = cgp_core_061 & input_e[0];
  assign cgp_core_065 = cgp_core_062 | cgp_core_064;
  assign cgp_core_066 = cgp_core_058 ^ cgp_core_065;
  assign cgp_core_067 = cgp_core_058 & cgp_core_065;
  assign cgp_core_068 = cgp_core_043 ^ cgp_core_059;
  assign cgp_core_069 = cgp_core_043 & cgp_core_059;
  assign cgp_core_070 = cgp_core_047 ^ cgp_core_063;
  assign cgp_core_071 = cgp_core_047 & cgp_core_063;
  assign cgp_core_072 = cgp_core_070 ^ cgp_core_069;
  assign cgp_core_073 = cgp_core_070 & cgp_core_069;
  assign cgp_core_074 = cgp_core_071 | cgp_core_073;
  assign cgp_core_075 = cgp_core_050 ^ cgp_core_066;
  assign cgp_core_076 = cgp_core_050 & cgp_core_066;
  assign cgp_core_077 = cgp_core_075 ^ cgp_core_074;
  assign cgp_core_078 = cgp_core_075 & cgp_core_074;
  assign cgp_core_079 = cgp_core_076 | cgp_core_078;
  assign cgp_core_080 = cgp_core_051 | cgp_core_067;
  assign cgp_core_081 = input_c[1] & cgp_core_067;
  assign cgp_core_082 = cgp_core_080 | cgp_core_079;
  assign cgp_core_083 = cgp_core_080 & input_a[1];
  assign cgp_core_084 = cgp_core_081 | cgp_core_083;
  assign cgp_core_086 = ~cgp_core_084;
  assign cgp_core_087 = ~cgp_core_082;
  assign cgp_core_088 = cgp_core_035 & cgp_core_087;
  assign cgp_core_090 = ~(cgp_core_035 ^ cgp_core_082);
  assign cgp_core_091 = cgp_core_090 & cgp_core_086;
  assign cgp_core_092 = ~cgp_core_077;
  assign cgp_core_093 = cgp_core_034 & cgp_core_092;
  assign cgp_core_094 = cgp_core_093 & cgp_core_091;
  assign cgp_core_095 = ~(cgp_core_034 ^ cgp_core_077);
  assign cgp_core_096 = cgp_core_095 & cgp_core_091;
  assign cgp_core_097 = ~cgp_core_072;
  assign cgp_core_098 = cgp_core_031 & cgp_core_097;
  assign cgp_core_099 = cgp_core_098 & cgp_core_096;
  assign cgp_core_100 = ~(cgp_core_031 ^ cgp_core_072);
  assign cgp_core_101 = cgp_core_100 & cgp_core_096;
  assign cgp_core_102 = ~(input_d[1] ^ input_d[1]);
  assign cgp_core_104 = cgp_core_027 & cgp_core_101;
  assign cgp_core_105_not = ~cgp_core_068;
  assign cgp_core_106 = cgp_core_105_not & cgp_core_101;
  assign cgp_core_107 = cgp_core_099 | cgp_core_094;
  assign cgp_core_108 = cgp_core_104 | cgp_core_107;
  assign cgp_core_109 = cgp_core_088 | cgp_core_106;
  assign cgp_core_110 = cgp_core_108 | cgp_core_109;

  assign cgp_out[0] = cgp_core_110;
endmodule