module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_036;
  wire cgp_core_038_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059_not;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081_not;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_095;

  assign cgp_core_018 = input_h[0] ^ input_c[0];
  assign cgp_core_019 = input_b[0] & input_c[0];
  assign cgp_core_020 = ~input_c[0];
  assign cgp_core_021 = ~(input_b[0] | input_b[1]);
  assign cgp_core_025 = input_h[1] ^ input_d[0];
  assign cgp_core_026 = ~(input_h[1] | input_c[0]);
  assign cgp_core_027 = input_a[1] ^ cgp_core_019;
  assign cgp_core_029 = cgp_core_027 | cgp_core_026;
  assign cgp_core_030 = ~(input_b[0] & input_h[1]);
  assign cgp_core_032 = ~(input_f[0] ^ input_g[1]);
  assign cgp_core_033 = input_g[0] & input_d[0];
  assign cgp_core_034_not = ~input_d[0];
  assign cgp_core_036 = input_f[0] ^ input_d[1];
  assign cgp_core_038_not = ~cgp_core_036;
  assign cgp_core_041 = input_f[1] ^ input_e[1];
  assign cgp_core_042 = input_d[0] & cgp_core_034_not;
  assign cgp_core_044 = input_d[1] & input_d[1];
  assign cgp_core_046 = input_d[0] & input_a[0];
  assign cgp_core_047 = ~(input_b[1] | input_g[1]);
  assign cgp_core_048 = input_f[1] ^ cgp_core_047;
  assign cgp_core_050 = ~(input_g[1] & input_f[0]);
  assign cgp_core_051 = ~(cgp_core_025 ^ input_e[1]);
  assign cgp_core_052 = cgp_core_029 | input_b[0];
  assign cgp_core_054 = ~(cgp_core_052 | input_d[0]);
  assign cgp_core_055 = input_h[0] & input_h[1];
  assign cgp_core_057 = cgp_core_032 ^ cgp_core_048;
  assign cgp_core_058 = input_c[0] & cgp_core_048;
  assign cgp_core_059_not = ~input_a[0];
  assign cgp_core_060 = input_g[0] & input_b[1];
  assign cgp_core_063 = input_c[1] & input_e[0];
  assign cgp_core_066 = input_d[1] | input_g[0];
  assign cgp_core_068 = input_e[0] & input_c[0];
  assign cgp_core_069 = input_a[1] ^ input_f[1];
  assign cgp_core_070 = input_e[1] & input_c[1];
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 | input_g[0];
  assign cgp_core_074 = ~cgp_core_066;
  assign cgp_core_077 = input_b[0] & cgp_core_074;
  assign cgp_core_079 = cgp_core_059_not & input_d[1];
  assign cgp_core_080 = cgp_core_079 & cgp_core_077;
  assign cgp_core_081_not = ~input_g[1];
  assign cgp_core_082 = ~(input_h[1] ^ cgp_core_077);
  assign cgp_core_083 = ~cgp_core_071;
  assign cgp_core_084 = input_d[0] & cgp_core_083;
  assign cgp_core_087 = input_e[1] ^ cgp_core_082;
  assign cgp_core_089 = cgp_core_050 & input_b[1];
  assign cgp_core_090 = input_g[1] | input_e[1];
  assign cgp_core_095 = ~(cgp_core_066 ^ input_g[0]);

  assign cgp_out[0] = 1'b1;
endmodule