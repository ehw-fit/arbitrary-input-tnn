module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_023_not;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031_not;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072_not;
  wire cgp_core_073;
  wire cgp_core_075;

  assign cgp_core_014 = ~input_a[5];
  assign cgp_core_015 = ~input_a[1];
  assign cgp_core_016 = input_a[9] | input_a[4];
  assign cgp_core_017 = ~(input_a[1] & input_a[7]);
  assign cgp_core_019 = ~(input_a[2] & input_a[4]);
  assign cgp_core_023_not = ~input_a[0];
  assign cgp_core_025 = input_a[6] | input_a[4];
  assign cgp_core_026 = ~(input_a[0] & input_a[5]);
  assign cgp_core_027 = ~input_a[2];
  assign cgp_core_028 = ~(input_a[0] ^ input_a[0]);
  assign cgp_core_029 = input_a[2] | input_a[9];
  assign cgp_core_030 = ~input_a[11];
  assign cgp_core_031_not = ~input_a[8];
  assign cgp_core_032 = input_a[4] | input_a[2];
  assign cgp_core_035 = ~(input_a[8] ^ input_a[11]);
  assign cgp_core_036 = input_a[5] ^ input_a[7];
  assign cgp_core_039 = ~input_a[6];
  assign cgp_core_040 = ~(input_a[2] ^ input_a[11]);
  assign cgp_core_041 = input_a[7] & input_a[6];
  assign cgp_core_042 = ~input_a[10];
  assign cgp_core_043 = ~(input_a[9] & input_a[7]);
  assign cgp_core_044 = ~input_a[10];
  assign cgp_core_045 = input_a[2] & input_a[4];
  assign cgp_core_046 = ~(input_a[8] ^ input_a[2]);
  assign cgp_core_047 = ~(input_a[0] & input_a[4]);
  assign cgp_core_049 = ~(input_a[9] ^ input_a[8]);
  assign cgp_core_051 = ~(input_a[3] ^ input_a[0]);
  assign cgp_core_052 = input_a[6] | input_a[2];
  assign cgp_core_053 = ~input_a[1];
  assign cgp_core_054 = input_a[8] & input_a[5];
  assign cgp_core_055 = ~(input_a[4] | input_a[1]);
  assign cgp_core_056 = input_a[10] | input_a[3];
  assign cgp_core_058 = input_a[11] | input_a[4];
  assign cgp_core_059 = input_a[7] ^ input_a[2];
  assign cgp_core_060 = ~input_a[11];
  assign cgp_core_064 = ~(input_a[4] | input_a[9]);
  assign cgp_core_065 = ~(input_a[9] ^ input_a[5]);
  assign cgp_core_068 = ~input_a[11];
  assign cgp_core_069 = input_a[8] & input_a[0];
  assign cgp_core_070 = input_a[5] ^ input_a[4];
  assign cgp_core_072_not = ~input_a[1];
  assign cgp_core_073 = input_a[2] & input_a[7];
  assign cgp_core_075 = ~(input_a[8] | input_a[6]);

  assign cgp_out[0] = 1'b1;
  assign cgp_out[1] = input_a[5];
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = 1'b0;
endmodule