module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_080;

  assign cgp_core_017 = input_a[0] ^ input_d[2];
  assign cgp_core_019 = input_a[1] | input_b[1];
  assign cgp_core_021 = ~(input_d[2] & input_a[2]);
  assign cgp_core_022 = ~(cgp_core_019 & input_e[1]);
  assign cgp_core_023 = input_a[1] & input_d[1];
  assign cgp_core_027 = input_b[1] & input_b[1];
  assign cgp_core_028 = input_a[2] | input_b[0];
  assign cgp_core_029 = input_d[0] ^ input_e[0];
  assign cgp_core_030 = input_c[2] & input_b[1];
  assign cgp_core_031 = input_d[1] & input_d[0];
  assign cgp_core_032 = input_c[2] | input_e[1];
  assign cgp_core_033 = input_c[1] ^ input_e[2];
  assign cgp_core_034 = ~(input_a[1] & cgp_core_030);
  assign cgp_core_035 = ~(input_e[0] & input_c[1]);
  assign cgp_core_036 = input_d[2] ^ input_d[0];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038 = cgp_core_036 ^ input_b[1];
  assign cgp_core_039 = input_e[0] ^ input_b[1];
  assign cgp_core_040 = input_b[0] | cgp_core_039;
  assign cgp_core_043 = input_c[1] ^ cgp_core_033;
  assign cgp_core_044 = input_c[1] & cgp_core_033;
  assign cgp_core_045 = cgp_core_043 & input_c[0];
  assign cgp_core_046 = cgp_core_043 & input_d[0];
  assign cgp_core_047 = input_b[1] | cgp_core_046;
  assign cgp_core_048 = input_c[2] ^ input_d[1];
  assign cgp_core_050 = cgp_core_048 ^ cgp_core_047;
  assign cgp_core_052 = ~(input_b[0] ^ input_a[1]);
  assign cgp_core_053 = ~cgp_core_040;
  assign cgp_core_054 = cgp_core_040 & input_a[1];
  assign cgp_core_055 = ~(input_a[2] | input_a[2]);
  assign cgp_core_057 = ~input_c[1];
  assign cgp_core_058 = cgp_core_028 & cgp_core_057;
  assign cgp_core_060 = ~(cgp_core_028 ^ input_d[2]);
  assign cgp_core_062 = cgp_core_050 ^ cgp_core_050;
  assign cgp_core_063 = input_e[0] & cgp_core_062;
  assign cgp_core_067 = ~(cgp_core_045 & input_a[1]);
  assign cgp_core_068 = cgp_core_021 | input_d[1];
  assign cgp_core_069 = ~input_d[0];
  assign cgp_core_070 = ~(cgp_core_021 ^ cgp_core_045);
  assign cgp_core_071 = input_b[1] ^ input_a[2];
  assign cgp_core_072 = ~input_d[1];
  assign cgp_core_073 = cgp_core_017 & cgp_core_072;
  assign cgp_core_074 = input_a[0] & input_e[0];
  assign cgp_core_075 = ~(input_c[0] & input_e[2]);
  assign cgp_core_080 = input_d[0] & input_c[0];

  assign cgp_out[0] = input_a[1];
endmodule