module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047_not;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055_not;

  assign cgp_core_014 = input_a[0] ^ input_a[0];
  assign cgp_core_015 = input_c[1] & input_b[2];
  assign cgp_core_016 = ~(input_a[2] | input_d[2]);
  assign cgp_core_018 = ~input_b[2];
  assign cgp_core_019 = ~input_c[2];
  assign cgp_core_020 = ~(input_c[2] & input_a[1]);
  assign cgp_core_021 = ~(input_d[2] | input_a[1]);
  assign cgp_core_023 = input_a[0] | input_a[2];
  assign cgp_core_025 = input_b[2] | input_a[2];
  assign cgp_core_026 = input_b[2] ^ input_d[1];
  assign cgp_core_027 = input_c[2] | input_a[0];
  assign cgp_core_032 = ~input_c[1];
  assign cgp_core_033 = input_c[2] | input_b[0];
  assign cgp_core_035 = ~input_b[2];
  assign cgp_core_036 = input_d[2] & input_c[2];
  assign cgp_core_038 = ~cgp_core_036;
  assign cgp_core_039 = cgp_core_025 & cgp_core_038;
  assign cgp_core_040 = ~(input_a[2] | input_b[2]);
  assign cgp_core_041 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_042_not = ~input_b[1];
  assign cgp_core_044 = ~(input_d[2] & input_c[0]);
  assign cgp_core_046 = input_a[0] & input_d[1];
  assign cgp_core_047_not = ~input_a[1];
  assign cgp_core_050 = ~input_d[1];
  assign cgp_core_052 = input_a[1] | input_a[1];
  assign cgp_core_054 = input_a[2] | input_a[2];
  assign cgp_core_055_not = ~input_c[2];

  assign cgp_out[0] = cgp_core_039;
endmodule