module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030_not;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_015 = input_b[1] & input_e[1];
  assign cgp_core_016 = input_d[1] & input_c[1];
  assign cgp_core_017 = input_a[1] & input_a[0];
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = input_a[1] & input_b[0];
  assign cgp_core_020 = input_d[1] & input_e[1];
  assign cgp_core_021 = ~(input_b[0] | input_e[1]);
  assign cgp_core_025 = input_c[0] & input_d[1];
  assign cgp_core_026 = ~(input_e[0] ^ input_b[1]);
  assign cgp_core_028 = ~input_c[0];
  assign cgp_core_030_not = ~input_c[0];
  assign cgp_core_032 = input_d[0] | input_d[0];
  assign cgp_core_034 = input_d[1] | input_c[1];
  assign cgp_core_035_not = ~input_b[1];
  assign cgp_core_036 = ~cgp_core_034;
  assign cgp_core_040 = input_c[1] & input_e[0];
  assign cgp_core_041 = input_c[1] | input_d[0];
  assign cgp_core_044 = input_b[1] | input_a[0];
  assign cgp_core_045 = ~input_e[1];
  assign cgp_core_053 = cgp_core_036 | cgp_core_018;
  assign cgp_core_054 = cgp_core_019 | cgp_core_053;

  assign cgp_out[0] = cgp_core_054;
endmodule