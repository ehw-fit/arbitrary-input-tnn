module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_018 = ~(input_b[2] | input_d[1]);
  assign cgp_core_020 = input_d[1] & input_a[1];
  assign cgp_core_021 = input_c[0] | input_e[2];
  assign cgp_core_022 = input_e[1] | input_e[2];
  assign cgp_core_023 = ~(input_d[0] & input_b[2]);
  assign cgp_core_024 = ~(input_a[0] | input_c[2]);
  assign cgp_core_025 = input_c[1] & input_c[0];
  assign cgp_core_026 = input_e[0] & input_b[2];
  assign cgp_core_027 = input_c[2] & input_b[2];
  assign cgp_core_028 = input_e[2] | cgp_core_027;
  assign cgp_core_029 = input_c[1] | input_c[2];
  assign cgp_core_030 = ~(input_d[1] ^ input_a[0]);
  assign cgp_core_032 = ~(input_b[0] | input_a[2]);
  assign cgp_core_035 = ~(input_e[2] & input_b[2]);
  assign cgp_core_038 = ~(input_b[0] ^ input_b[0]);
  assign cgp_core_039 = ~(input_c[0] ^ input_a[2]);
  assign cgp_core_040 = ~(input_d[0] | input_c[0]);
  assign cgp_core_041 = input_b[2] | input_c[2];
  assign cgp_core_043 = ~input_d[1];
  assign cgp_core_044 = ~(input_a[1] & input_e[2]);
  assign cgp_core_045 = input_a[1] | input_a[0];
  assign cgp_core_047 = ~input_a[2];
  assign cgp_core_048_not = ~input_a[0];
  assign cgp_core_049 = input_c[1] ^ input_b[2];
  assign cgp_core_050 = ~input_a[0];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_056 = ~cgp_core_051;
  assign cgp_core_057 = cgp_core_041 & cgp_core_056;
  assign cgp_core_059 = ~(input_c[1] | input_c[1]);
  assign cgp_core_060 = input_b[2] & input_c[2];
  assign cgp_core_064 = ~(input_c[0] | input_e[1]);
  assign cgp_core_067 = input_b[0] & input_d[1];
  assign cgp_core_069_not = ~input_e[0];
  assign cgp_core_070 = ~(input_a[0] ^ input_b[2]);
  assign cgp_core_071 = ~input_c[1];
  assign cgp_core_072 = ~(input_b[0] | input_d[2]);
  assign cgp_core_073 = ~(input_c[1] | input_e[1]);
  assign cgp_core_076 = ~(input_b[0] & input_b[1]);
  assign cgp_core_079 = cgp_core_057 | cgp_core_028;
  assign cgp_core_080 = ~(input_d[2] | input_e[2]);

  assign cgp_out[0] = cgp_core_079;
endmodule