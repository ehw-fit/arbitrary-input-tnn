module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_031_not;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_044_not;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;
  wire cgp_core_097;

  assign cgp_core_021 = input_c[0] | input_f[1];
  assign cgp_core_022 = input_e[0] | input_c[1];
  assign cgp_core_024 = ~(input_e[0] ^ input_e[0]);
  assign cgp_core_025 = ~input_a[2];
  assign cgp_core_027 = ~(input_f[2] | input_b[0]);
  assign cgp_core_029 = input_b[2] & input_d[0];
  assign cgp_core_031_not = ~input_e[2];
  assign cgp_core_033 = ~(input_f[2] | input_d[1]);
  assign cgp_core_034 = input_b[2] | input_e[2];
  assign cgp_core_036 = ~input_e[2];
  assign cgp_core_037_not = ~input_b[0];
  assign cgp_core_039 = input_b[2] | input_f[0];
  assign cgp_core_042 = ~(input_d[1] & input_b[2]);
  assign cgp_core_044_not = ~input_b[2];
  assign cgp_core_046 = ~input_a[0];
  assign cgp_core_047 = ~(input_b[1] | input_d[1]);
  assign cgp_core_048 = input_e[2] ^ input_a[1];
  assign cgp_core_049 = input_e[1] ^ input_f[2];
  assign cgp_core_053 = input_c[0] & input_b[1];
  assign cgp_core_055 = input_a[0] | input_b[0];
  assign cgp_core_056 = ~(input_f[1] & input_c[1]);
  assign cgp_core_057 = input_a[1] ^ input_f[0];
  assign cgp_core_058 = ~(input_e[1] & input_e[0]);
  assign cgp_core_060 = ~input_f[0];
  assign cgp_core_062 = ~input_e[2];
  assign cgp_core_064 = ~(input_a[2] | input_e[2]);
  assign cgp_core_071 = ~(input_a[1] ^ input_d[2]);
  assign cgp_core_072 = ~(input_e[2] ^ input_a[2]);
  assign cgp_core_074 = input_f[0] ^ input_c[2];
  assign cgp_core_075 = ~(input_a[0] ^ input_b[1]);
  assign cgp_core_077 = input_e[0] ^ input_d[1];
  assign cgp_core_078 = ~input_c[2];
  assign cgp_core_079 = ~input_f[1];
  assign cgp_core_080 = ~input_d[2];
  assign cgp_core_081 = ~(input_b[1] & input_b[0]);
  assign cgp_core_082 = input_a[1] & input_e[0];
  assign cgp_core_083 = ~(input_d[2] ^ input_c[1]);
  assign cgp_core_084 = ~input_c[1];
  assign cgp_core_085 = ~(input_a[2] | input_d[2]);
  assign cgp_core_088 = input_d[2] | input_e[0];
  assign cgp_core_090 = input_a[1] & input_b[1];
  assign cgp_core_091 = ~input_a[0];
  assign cgp_core_093 = input_a[2] & input_a[2];
  assign cgp_core_097 = ~(input_c[2] ^ input_d[0]);

  assign cgp_out[0] = input_a[1];
endmodule