module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035_not;
  wire cgp_core_037_not;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046_not;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;

  assign cgp_core_014 = input_b[1] ^ input_f[0];
  assign cgp_core_015 = input_b[1] & input_a[0];
  assign cgp_core_016 = input_b[0] ^ input_a[0];
  assign cgp_core_018 = cgp_core_016 ^ cgp_core_015;
  assign cgp_core_019 = cgp_core_016 & cgp_core_015;
  assign cgp_core_021 = input_e[0] | input_b[0];
  assign cgp_core_022 = input_e[0] & input_f[0];
  assign cgp_core_024 = input_e[1] & input_b[0];
  assign cgp_core_025 = input_d[0] ^ cgp_core_022;
  assign cgp_core_026 = input_e[1] & cgp_core_022;
  assign cgp_core_027 = cgp_core_024 | cgp_core_026;
  assign cgp_core_029 = input_d[0] & input_f[0];
  assign cgp_core_030 = input_d[1] ^ cgp_core_025;
  assign cgp_core_031 = ~(input_d[1] | cgp_core_025);
  assign cgp_core_032 = cgp_core_030 ^ cgp_core_029;
  assign cgp_core_033 = cgp_core_030 & cgp_core_029;
  assign cgp_core_035_not = ~cgp_core_027;
  assign cgp_core_037_not = ~cgp_core_014;
  assign cgp_core_039 = ~input_a[0];
  assign cgp_core_040 = cgp_core_018 & cgp_core_032;
  assign cgp_core_041 = cgp_core_039 ^ input_e[0];
  assign cgp_core_044 = cgp_core_019 & cgp_core_035_not;
  assign cgp_core_045 = cgp_core_019 & cgp_core_035_not;
  assign cgp_core_046_not = ~cgp_core_044;
  assign cgp_core_047 = cgp_core_044 & input_e[0];
  assign cgp_core_051 = ~input_d[1];
  assign cgp_core_056 = ~(cgp_core_046_not | cgp_core_046_not);
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_061 = ~(cgp_core_041 ^ input_b[1]);
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_064 = cgp_core_037_not & input_e[1];
  assign cgp_core_065 = cgp_core_064 & input_a[1];
  assign cgp_core_066 = ~(cgp_core_037_not ^ input_e[1]);
  assign cgp_core_067 = cgp_core_066 & input_f[0];
  assign cgp_core_068 = input_f[1] | cgp_core_046_not;

  assign cgp_out[0] = 1'b1;
endmodule