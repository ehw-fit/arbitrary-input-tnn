module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_080_not;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_096;
  wire cgp_core_098;
  wire cgp_core_103;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_108;
  wire cgp_core_110;

  assign cgp_core_021 = input_h[0] & input_i[0];
  assign cgp_core_023 = ~(input_f[0] & input_a[1]);
  assign cgp_core_027 = input_d[0] ^ input_i[1];
  assign cgp_core_029 = ~(input_d[1] & input_i[1]);
  assign cgp_core_030 = ~input_d[1];
  assign cgp_core_032 = input_b[0] & input_d[0];
  assign cgp_core_033 = cgp_core_030 | cgp_core_032;
  assign cgp_core_036 = input_b[0] ^ input_a[1];
  assign cgp_core_037 = input_b[0] & input_c[1];
  assign cgp_core_038 = ~input_g[0];
  assign cgp_core_039 = ~(input_h[0] & input_c[0]);
  assign cgp_core_041 = ~input_a[0];
  assign cgp_core_042 = ~(cgp_core_039 ^ cgp_core_041);
  assign cgp_core_043 = input_g[0] & input_d[1];
  assign cgp_core_044 = input_g[0] & input_e[1];
  assign cgp_core_045_not = ~input_c[0];
  assign cgp_core_046 = ~(input_c[1] & input_f[1]);
  assign cgp_core_048 = ~(input_c[0] ^ cgp_core_044);
  assign cgp_core_049 = input_b[1] & input_f[0];
  assign cgp_core_050 = ~(input_b[0] | cgp_core_049);
  assign cgp_core_051 = input_b[1] & input_f[1];
  assign cgp_core_053 = ~(input_f[1] ^ input_f[0]);
  assign cgp_core_054 = ~(input_e[0] ^ input_c[0]);
  assign cgp_core_055 = input_f[1] | input_b[1];
  assign cgp_core_057 = input_a[0] | input_e[0];
  assign cgp_core_058 = input_b[1] | input_g[0];
  assign cgp_core_060 = input_i[0] & input_e[1];
  assign cgp_core_061 = input_b[1] | input_e[0];
  assign cgp_core_062 = ~input_g[0];
  assign cgp_core_063 = input_a[1] ^ input_i[1];
  assign cgp_core_064 = ~input_b[1];
  assign cgp_core_066 = input_g[1] ^ input_e[0];
  assign cgp_core_068 = ~(cgp_core_043 | input_c[0]);
  assign cgp_core_070 = input_c[1] ^ cgp_core_063;
  assign cgp_core_071 = input_a[1] & input_f[1];
  assign cgp_core_072 = ~cgp_core_070;
  assign cgp_core_073 = ~(input_g[1] | input_b[0]);
  assign cgp_core_076 = ~(input_b[0] & input_f[0]);
  assign cgp_core_080_not = ~input_h[0];
  assign cgp_core_082 = ~input_f[1];
  assign cgp_core_083 = input_h[1] & input_f[0];
  assign cgp_core_084 = input_d[0] | input_c[1];
  assign cgp_core_085 = ~(cgp_core_084 ^ input_i[0]);
  assign cgp_core_086 = ~input_a[0];
  assign cgp_core_087 = ~(input_h[1] | input_b[1]);
  assign cgp_core_089 = input_b[0] & input_a[0];
  assign cgp_core_090 = ~(input_b[0] ^ input_f[1]);
  assign cgp_core_091 = input_b[1] & input_h[1];
  assign cgp_core_092 = ~(input_i[0] | input_c[0]);
  assign cgp_core_096 = input_h[0] & input_c[0];
  assign cgp_core_098 = ~input_c[0];
  assign cgp_core_103 = ~input_c[0];
  assign cgp_core_104 = input_g[1] & input_h[1];
  assign cgp_core_105 = ~(cgp_core_027 | input_c[1]);
  assign cgp_core_106 = ~input_h[0];
  assign cgp_core_108 = input_i[0] | input_i[0];
  assign cgp_core_110 = ~(input_h[1] & input_g[0]);

  assign cgp_out[0] = 1'b0;
endmodule