module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_016 = ~(input_d[1] & input_d[2]);
  assign cgp_core_017 = input_d[1] ^ input_b[1];
  assign cgp_core_019 = input_a[0] | input_d[1];
  assign cgp_core_023 = ~input_c[2];
  assign cgp_core_024 = ~(input_c[1] & input_a[2]);
  assign cgp_core_026 = ~(input_b[0] | input_d[0]);
  assign cgp_core_027 = ~(input_b[2] | input_c[2]);
  assign cgp_core_030 = ~(input_d[0] | input_d[2]);
  assign cgp_core_033 = ~(input_d[1] ^ input_c[0]);
  assign cgp_core_034 = ~input_c[1];
  assign cgp_core_035 = input_b[2] | input_b[0];
  assign cgp_core_038 = input_d[2] | input_b[1];
  assign cgp_core_041 = ~(input_c[0] & input_d[1]);
  assign cgp_core_044 = ~(input_a[1] | input_b[1]);
  assign cgp_core_046 = input_b[0] & input_d[2];
  assign cgp_core_047 = input_b[1] & input_c[2];
  assign cgp_core_048 = ~input_c[2];
  assign cgp_core_049 = input_a[1] | input_a[1];
  assign cgp_core_050 = input_b[1] & input_d[2];
  assign cgp_core_052 = ~(input_d[1] & input_a[2]);
  assign cgp_core_055 = ~input_a[0];
  assign cgp_core_056 = ~(input_a[2] | input_c[1]);
  assign cgp_core_058 = input_d[2] & input_b[2];
  assign cgp_core_059 = ~(input_a[1] | input_d[2]);

  assign cgp_out[0] = input_b[2];
endmodule