module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;

  assign cgp_core_011 = input_c[0] & input_d[0];
  assign cgp_core_012 = input_c[1] | input_d[1];
  assign cgp_core_013 = input_c[1] & input_d[1];
  assign cgp_core_014 = cgp_core_012 | cgp_core_011;
  assign cgp_core_015 = cgp_core_012 & input_d[0];
  assign cgp_core_016 = cgp_core_013 | cgp_core_015;
  assign cgp_core_018 = input_b[0] & input_a[0];
  assign cgp_core_019 = input_b[1] | cgp_core_014;
  assign cgp_core_020 = input_b[1] & cgp_core_014;
  assign cgp_core_021 = cgp_core_019 | cgp_core_018;
  assign cgp_core_022 = cgp_core_019 & input_b[0];
  assign cgp_core_023 = cgp_core_020 | cgp_core_022;
  assign cgp_core_024 = cgp_core_016 | cgp_core_023;
  assign cgp_core_026 = input_b[0] | input_d[1];
  assign cgp_core_030 = ~input_a[1];
  assign cgp_core_031 = cgp_core_021 & cgp_core_030;
  assign cgp_core_033 = ~(cgp_core_021 ^ input_a[1]);
  assign cgp_core_035 = ~input_a[0];
  assign cgp_core_037 = cgp_core_035 & cgp_core_033;
  assign cgp_core_039 = ~(input_d[0] & input_b[0]);
  assign cgp_core_040 = cgp_core_037 | cgp_core_031;
  assign cgp_core_041 = input_a[1] | input_d[1];
  assign cgp_core_043 = cgp_core_040 | cgp_core_024;

  assign cgp_out[0] = cgp_core_043;
endmodule