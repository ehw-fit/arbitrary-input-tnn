module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038_not;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_073;
  wire cgp_core_076;

  assign cgp_core_017 = input_b[0] ^ input_d[0];
  assign cgp_core_018 = input_b[0] & input_c[0];
  assign cgp_core_019 = input_b[2] ^ input_c[1];
  assign cgp_core_021 = cgp_core_019 ^ input_d[2];
  assign cgp_core_022 = cgp_core_019 & input_e[0];
  assign cgp_core_023 = input_b[2] | input_a[2];
  assign cgp_core_024 = input_a[1] ^ input_c[2];
  assign cgp_core_025 = input_b[2] & input_c[0];
  assign cgp_core_027 = cgp_core_024 ^ input_e[1];
  assign cgp_core_029 = ~input_d[0];
  assign cgp_core_030 = ~(input_c[1] | input_e[0]);
  assign cgp_core_031 = input_d[1] | input_e[1];
  assign cgp_core_032 = input_c[2] & input_e[1];
  assign cgp_core_033 = ~cgp_core_031;
  assign cgp_core_034 = ~(input_e[2] | input_a[0]);
  assign cgp_core_035 = ~cgp_core_032;
  assign cgp_core_036 = input_e[0] ^ input_a[2];
  assign cgp_core_037 = input_e[0] & input_e[2];
  assign cgp_core_038_not = ~cgp_core_036;
  assign cgp_core_039 = cgp_core_036 & input_b[1];
  assign cgp_core_040 = ~(cgp_core_037 & cgp_core_039);
  assign cgp_core_041 = input_e[2] ^ input_a[2];
  assign cgp_core_042 = cgp_core_017 & cgp_core_029;
  assign cgp_core_043_not = ~cgp_core_033;
  assign cgp_core_044 = cgp_core_021 & cgp_core_033;
  assign cgp_core_045 = ~input_c[0];
  assign cgp_core_046 = cgp_core_043_not & input_d[1];
  assign cgp_core_048 = ~(cgp_core_023 | cgp_core_038_not);
  assign cgp_core_049 = cgp_core_023 & cgp_core_038_not;
  assign cgp_core_050_not = ~cgp_core_048;
  assign cgp_core_066 = input_c[0] ^ cgp_core_050_not;
  assign cgp_core_068 = ~(cgp_core_045 | cgp_core_045);
  assign cgp_core_073 = ~cgp_core_041;
  assign cgp_core_076 = ~input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule