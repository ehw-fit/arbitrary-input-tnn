module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039_not;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[0] ^ input_a[9];
  assign cgp_core_020 = ~(input_a[7] | input_a[5]);
  assign cgp_core_021 = ~(input_a[8] ^ input_a[5]);
  assign cgp_core_023 = input_a[11] ^ input_a[0];
  assign cgp_core_026 = ~input_a[7];
  assign cgp_core_027 = ~(input_a[4] ^ input_a[2]);
  assign cgp_core_028 = ~input_a[0];
  assign cgp_core_031 = ~(input_a[6] & input_a[10]);
  assign cgp_core_032 = ~(input_a[11] & input_a[11]);
  assign cgp_core_033 = input_a[8] ^ input_a[3];
  assign cgp_core_034 = ~(input_a[7] | input_a[9]);
  assign cgp_core_036 = ~(input_a[2] & input_a[0]);
  assign cgp_core_038 = ~(input_a[0] & input_a[5]);
  assign cgp_core_039_not = ~input_a[6];
  assign cgp_core_040 = ~input_a[3];
  assign cgp_core_042 = ~(input_a[11] ^ input_a[3]);
  assign cgp_core_044 = ~(input_a[4] & input_a[4]);
  assign cgp_core_047 = input_a[8] | input_a[10];
  assign cgp_core_051 = ~(input_a[11] | input_a[0]);
  assign cgp_core_052 = ~(input_a[7] & input_a[2]);
  assign cgp_core_053 = input_a[3] ^ input_a[3];
  assign cgp_core_058 = ~(input_a[8] & input_a[6]);
  assign cgp_core_059 = input_a[10] ^ input_a[6];
  assign cgp_core_060 = ~input_a[8];
  assign cgp_core_062 = input_a[0] & input_a[1];
  assign cgp_core_063 = ~(input_a[4] & input_a[6]);
  assign cgp_core_065 = input_a[6] ^ input_a[6];
  assign cgp_core_066 = ~input_a[10];
  assign cgp_core_068 = input_a[10] & input_a[8];
  assign cgp_core_073 = input_a[5] ^ input_a[2];
  assign cgp_core_074 = input_a[4] | input_a[11];
  assign cgp_core_077 = ~(input_a[1] & input_a[4]);
  assign cgp_core_078 = ~(input_a[9] ^ input_a[5]);

  assign cgp_out[0] = 1'b1;
  assign cgp_out[1] = 1'b1;
  assign cgp_out[2] = input_a[0];
  assign cgp_out[3] = 1'b0;
endmodule