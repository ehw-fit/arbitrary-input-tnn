module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_025 = ~(input_a[4] & input_a[3]);
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_037 = input_a[7] & input_a[0];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_043 = ~input_a[5];
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_060 = input_a[11] & input_a[9];
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~(input_a[9] ^ input_a[5]);
  assign cgp_core_075 = ~input_a[1];
  assign cgp_core_076 = ~(input_a[3] ^ input_a[8]);
  assign cgp_core_078 = ~(input_a[5] | input_a[8]);

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule