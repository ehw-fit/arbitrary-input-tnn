module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_037_not;
  wire cgp_core_038;
  wire cgp_core_039_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058_not;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_083;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_021 = input_e[1] ^ input_d[2];
  assign cgp_core_025 = ~(input_e[0] | input_b[2]);
  assign cgp_core_027 = input_c[2] | input_e[2];
  assign cgp_core_028 = input_c[2] & input_e[2];
  assign cgp_core_029 = ~(input_c[2] | input_d[2]);
  assign cgp_core_030 = cgp_core_027 & input_a[2];
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = input_c[1] & input_c[2];
  assign cgp_core_037_not = ~input_b[2];
  assign cgp_core_038 = ~(input_e[2] | input_b[2]);
  assign cgp_core_039_not = ~input_b[0];
  assign cgp_core_041 = input_d[1] ^ input_f[0];
  assign cgp_core_042 = ~(input_c[1] | input_f[2]);
  assign cgp_core_043 = ~(input_d[1] & input_d[0]);
  assign cgp_core_047 = ~input_c[1];
  assign cgp_core_048 = input_c[0] | input_f[1];
  assign cgp_core_049 = input_d[1] & input_e[0];
  assign cgp_core_050 = input_d[1] & input_b[2];
  assign cgp_core_051 = ~input_a[1];
  assign cgp_core_052 = ~(input_f[2] | input_f[0]);
  assign cgp_core_053 = input_d[2] | input_f[2];
  assign cgp_core_054 = input_d[2] & input_f[2];
  assign cgp_core_056 = cgp_core_053 & input_f[1];
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058_not = ~input_e[2];
  assign cgp_core_059 = input_a[0] ^ input_d[0];
  assign cgp_core_060 = input_e[2] & input_b[0];
  assign cgp_core_061 = ~(input_f[1] | input_b[1]);
  assign cgp_core_062 = input_e[0] | input_f[1];
  assign cgp_core_065 = ~(input_d[1] ^ input_f[1]);
  assign cgp_core_067 = ~(input_d[0] ^ input_d[0]);
  assign cgp_core_068 = ~(input_c[2] ^ input_e[2]);
  assign cgp_core_069 = input_c[2] | input_b[2];
  assign cgp_core_070 = cgp_core_057 | input_b[2];
  assign cgp_core_071 = cgp_core_057 & input_b[2];
  assign cgp_core_072 = ~cgp_core_071;
  assign cgp_core_073 = cgp_core_031 & cgp_core_072;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_078 = ~(input_b[1] & input_d[0]);
  assign cgp_core_083 = input_a[1] ^ input_a[0];
  assign cgp_core_087 = ~(input_f[0] & input_f[1]);
  assign cgp_core_088 = input_b[1] & input_f[0];
  assign cgp_core_089 = ~(input_f[0] & input_a[1]);
  assign cgp_core_090 = ~input_e[0];
  assign cgp_core_091 = input_a[0] | input_d[1];
  assign cgp_core_093 = ~(input_c[1] ^ input_d[1]);
  assign cgp_core_095 = ~input_a[1];
  assign cgp_core_096 = ~(input_b[1] & input_f[2]);
  assign cgp_core_098 = cgp_core_075 | cgp_core_073;
  assign cgp_core_099 = input_d[2] & input_d[1];

  assign cgp_out[0] = cgp_core_098;
endmodule