module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_071_not;
  wire cgp_core_072_not;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;

  assign cgp_core_018 = ~(input_a[1] & input_a[0]);
  assign cgp_core_021 = ~input_b[0];
  assign cgp_core_023 = input_a[0] | input_a[1];
  assign cgp_core_026 = input_a[1] & input_d[1];
  assign cgp_core_027 = ~(input_d[0] | input_d[1]);
  assign cgp_core_031 = input_e[1] & cgp_core_026;
  assign cgp_core_032 = ~(input_c[0] | input_d[0]);
  assign cgp_core_033 = ~(input_c[0] ^ input_g[1]);
  assign cgp_core_034 = input_d[1] & input_f[1];
  assign cgp_core_035 = input_g[0] ^ input_e[1];
  assign cgp_core_036 = ~(input_c[0] | input_g[1]);
  assign cgp_core_037 = input_e[1] | input_d[1];
  assign cgp_core_039 = ~input_c[0];
  assign cgp_core_041 = ~(input_d[0] & input_d[0]);
  assign cgp_core_042_not = ~input_e[0];
  assign cgp_core_043 = ~(input_d[1] ^ input_c[0]);
  assign cgp_core_044 = input_g[1] ^ input_f[0];
  assign cgp_core_047 = input_b[0] | input_e[0];
  assign cgp_core_048 = ~(input_a[1] & input_c[0]);
  assign cgp_core_052 = input_b[1] ^ input_g[0];
  assign cgp_core_054 = input_e[0] | input_a[1];
  assign cgp_core_055 = input_c[0] & input_c[0];
  assign cgp_core_058 = ~(input_g[0] & input_g[0]);
  assign cgp_core_060 = ~(input_e[1] ^ input_f[1]);
  assign cgp_core_061 = ~input_a[0];
  assign cgp_core_062 = ~(input_b[0] | input_c[1]);
  assign cgp_core_064_not = ~input_c[0];
  assign cgp_core_065 = ~(input_b[0] & input_e[0]);
  assign cgp_core_066 = input_f[0] & input_e[1];
  assign cgp_core_068 = input_c[1] | input_d[1];
  assign cgp_core_071_not = ~input_e[1];
  assign cgp_core_072_not = ~input_d[1];
  assign cgp_core_074 = ~(input_d[0] ^ input_a[0]);
  assign cgp_core_075 = ~(input_d[0] | input_c[0]);
  assign cgp_core_078 = ~(input_c[0] & input_f[1]);

  assign cgp_out[0] = cgp_core_031;
endmodule