module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_051_not;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;

  assign cgp_core_017 = input_g[1] | input_c[0];
  assign cgp_core_018 = input_a[1] ^ input_g[0];
  assign cgp_core_020 = ~(cgp_core_018 | input_d[1]);
  assign cgp_core_021 = cgp_core_018 & input_g[1];
  assign cgp_core_022 = input_a[1] | input_c[0];
  assign cgp_core_023 = input_e[0] ^ input_b[1];
  assign cgp_core_026 = input_a[0] & input_g[1];
  assign cgp_core_027 = ~(input_a[1] ^ input_e[1]);
  assign cgp_core_030 = input_d[0] ^ cgp_core_023;
  assign cgp_core_031 = input_f[1] & cgp_core_023;
  assign cgp_core_032 = ~(input_g[0] ^ cgp_core_027);
  assign cgp_core_033 = input_d[1] & cgp_core_027;
  assign cgp_core_034 = cgp_core_032 ^ cgp_core_031;
  assign cgp_core_035 = cgp_core_032 & input_e[1];
  assign cgp_core_036 = cgp_core_033 | cgp_core_035;
  assign cgp_core_037 = ~(input_b[1] & cgp_core_036);
  assign cgp_core_038 = input_f[0] | cgp_core_036;
  assign cgp_core_039 = ~input_b[0];
  assign cgp_core_040 = input_b[1] & input_b[0];
  assign cgp_core_041 = ~(input_f[0] ^ cgp_core_034);
  assign cgp_core_042 = ~(cgp_core_020 & cgp_core_034);
  assign cgp_core_043 = input_e[0] ^ cgp_core_040;
  assign cgp_core_045 = input_c[0] | input_e[0];
  assign cgp_core_049 = input_f[0] & cgp_core_045;
  assign cgp_core_051_not = ~input_b[0];
  assign cgp_core_055 = input_f[0] ^ input_f[0];
  assign cgp_core_056 = ~(input_b[1] ^ input_f[1]);
  assign cgp_core_057 = input_c[1] ^ input_g[1];
  assign cgp_core_058 = cgp_core_055 & input_a[1];
  assign cgp_core_059 = input_g[1] | cgp_core_058;
  assign cgp_core_060 = ~cgp_core_038;
  assign cgp_core_061 = input_g[0] & cgp_core_060;
  assign cgp_core_062 = input_b[0] ^ cgp_core_051_not;
  assign cgp_core_063 = cgp_core_062 | cgp_core_060;
  assign cgp_core_064 = ~cgp_core_059;
  assign cgp_core_065 = input_c[1] & cgp_core_064;
  assign cgp_core_066 = cgp_core_065 & cgp_core_063;
  assign cgp_core_069 = ~input_a[0];
  assign cgp_core_070 = ~(input_d[0] | cgp_core_069);
  assign cgp_core_071 = input_g[0] & input_a[1];
  assign cgp_core_072 = ~(input_g[1] ^ input_e[1]);
  assign cgp_core_073 = cgp_core_072 & input_e[1];
  assign cgp_core_075 = ~cgp_core_039;
  assign cgp_core_076 = input_e[0] & cgp_core_073;
  assign cgp_core_077 = ~cgp_core_039;
  assign cgp_core_078 = cgp_core_077 & cgp_core_073;
  assign cgp_core_079 = ~cgp_core_071;
  assign cgp_core_080 = ~(input_b[1] | input_f[1]);
  assign cgp_core_081 = cgp_core_038 | input_b[1];

  assign cgp_out[0] = 1'b1;
endmodule