module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060_not;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = ~(input_a[1] ^ input_e[0]);
  assign cgp_core_018 = input_c[1] ^ input_d[1];
  assign cgp_core_019 = input_c[1] & input_d[1];
  assign cgp_core_020 = cgp_core_018 ^ input_g[1];
  assign cgp_core_021 = cgp_core_018 & input_g[1];
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_024 = input_e[1] | input_a[1];
  assign cgp_core_029 = input_a[1] ^ input_e[0];
  assign cgp_core_031 = ~(input_a[1] | input_a[0]);
  assign cgp_core_032 = ~cgp_core_020;
  assign cgp_core_034 = ~(cgp_core_032 & input_e[1]);
  assign cgp_core_035 = ~(input_b[1] & input_g[1]);
  assign cgp_core_036 = cgp_core_020 | input_e[1];
  assign cgp_core_039 = cgp_core_022 | input_e[1];
  assign cgp_core_040 = cgp_core_022 & cgp_core_036;
  assign cgp_core_043 = input_b[0] & input_a[0];
  assign cgp_core_044 = input_b[1] ^ input_f[1];
  assign cgp_core_045 = input_b[1] & input_f[1];
  assign cgp_core_046 = cgp_core_044 ^ cgp_core_043;
  assign cgp_core_047 = cgp_core_044 & cgp_core_043;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_049 = ~(input_d[0] | input_e[0]);
  assign cgp_core_050 = input_d[0] ^ input_g[0];
  assign cgp_core_051 = input_a[1] ^ cgp_core_046;
  assign cgp_core_052 = input_a[1] & cgp_core_046;
  assign cgp_core_054_not = ~input_g[0];
  assign cgp_core_056 = cgp_core_048 ^ cgp_core_052;
  assign cgp_core_057 = input_a[1] & input_f[1];
  assign cgp_core_060_not = ~cgp_core_057;
  assign cgp_core_061 = ~cgp_core_056;
  assign cgp_core_063 = cgp_core_061 & cgp_core_060_not;
  assign cgp_core_064 = cgp_core_039 & cgp_core_056;
  assign cgp_core_066 = ~cgp_core_051;
  assign cgp_core_067 = cgp_core_034 & cgp_core_066;
  assign cgp_core_068 = cgp_core_067 & cgp_core_064;
  assign cgp_core_069 = ~(input_a[0] ^ input_d[0]);
  assign cgp_core_072 = input_c[0] ^ input_b[1];
  assign cgp_core_074 = input_b[0] & input_a[0];
  assign cgp_core_078 = cgp_core_063 | cgp_core_040;
  assign cgp_core_079 = cgp_core_068 | cgp_core_078;

  assign cgp_out[0] = cgp_core_079;
endmodule