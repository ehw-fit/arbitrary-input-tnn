module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033_not;
  wire cgp_core_036;
  wire cgp_core_038_not;
  wire cgp_core_039;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_012 = input_d[1] ^ input_c[0];
  assign cgp_core_014 = input_b[0] | input_d[1];
  assign cgp_core_015 = input_a[0] & input_e[0];
  assign cgp_core_016 = ~(input_d[1] & input_b[0]);
  assign cgp_core_019 = input_c[0] ^ input_e[0];
  assign cgp_core_020 = input_c[0] | input_b[0];
  assign cgp_core_021 = input_c[1] ^ input_e[0];
  assign cgp_core_023 = ~(input_d[1] ^ input_e[0]);
  assign cgp_core_024 = cgp_core_021 & input_b[0];
  assign cgp_core_029 = input_a[1] & cgp_core_023;
  assign cgp_core_031 = ~input_e[0];
  assign cgp_core_033_not = ~input_a[1];
  assign cgp_core_036 = ~input_c[1];
  assign cgp_core_038_not = ~input_a[1];
  assign cgp_core_039 = cgp_core_038_not & input_d[0];
  assign cgp_core_043 = input_d[0] | input_a[0];
  assign cgp_core_046 = ~(cgp_core_016 ^ input_c[0]);
  assign cgp_core_048 = ~(input_c[0] | input_d[1]);
  assign cgp_core_052 = cgp_core_048 | input_b[1];
  assign cgp_core_053 = ~(cgp_core_039 ^ input_b[0]);
  assign cgp_core_054 = ~(input_a[0] ^ input_d[0]);

  assign cgp_out[0] = input_d[0];
endmodule