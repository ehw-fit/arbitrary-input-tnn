module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020_not;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_034;
  wire cgp_core_036_not;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_080;
  wire cgp_core_085;
  wire cgp_core_090;
  wire cgp_core_091;

  assign cgp_core_020_not = ~input_b[0];
  assign cgp_core_023 = input_b[0] & input_e[2];
  assign cgp_core_025 = ~(input_a[1] | input_c[0]);
  assign cgp_core_027 = ~(input_d[0] | input_c[0]);
  assign cgp_core_028 = input_a[2] & input_b[2];
  assign cgp_core_034 = input_a[0] | input_e[1];
  assign cgp_core_036_not = ~cgp_core_034;
  assign cgp_core_037 = ~(cgp_core_034 | input_c[0]);
  assign cgp_core_039 = input_f[2] & input_d[2];
  assign cgp_core_040 = input_a[0] & input_f[2];
  assign cgp_core_042 = input_e[1] ^ input_b[1];
  assign cgp_core_043 = input_e[1] | input_d[1];
  assign cgp_core_045 = ~(input_b[1] ^ input_e[0]);
  assign cgp_core_046 = input_d[0] | input_a[0];
  assign cgp_core_047 = ~input_e[1];
  assign cgp_core_049 = input_b[1] & cgp_core_045;
  assign cgp_core_050 = cgp_core_047 | cgp_core_049;
  assign cgp_core_051 = input_a[1] & input_f[0];
  assign cgp_core_052 = ~(input_e[2] ^ input_a[0]);
  assign cgp_core_053 = ~(input_e[2] ^ cgp_core_050);
  assign cgp_core_054 = input_a[2] & cgp_core_050;
  assign cgp_core_055 = input_b[1] | input_a[0];
  assign cgp_core_057 = input_a[2] & input_e[1];
  assign cgp_core_058 = input_d[0] ^ input_a[2];
  assign cgp_core_059 = cgp_core_036_not ^ input_a[0];
  assign cgp_core_060 = ~(input_a[0] | cgp_core_057);
  assign cgp_core_061 = cgp_core_058 ^ cgp_core_057;
  assign cgp_core_064 = ~input_b[1];
  assign cgp_core_067 = ~(input_c[1] | input_e[1]);
  assign cgp_core_068 = cgp_core_043 | input_a[2];
  assign cgp_core_069 = input_d[1] & input_d[0];
  assign cgp_core_070 = cgp_core_068 ^ input_d[2];
  assign cgp_core_071 = ~(cgp_core_068 & input_e[0]);
  assign cgp_core_073 = ~input_a[2];
  assign cgp_core_075 = ~input_b[2];
  assign cgp_core_080 = ~input_f[1];
  assign cgp_core_085 = ~input_c[1];
  assign cgp_core_090 = ~(input_e[0] | input_f[2]);
  assign cgp_core_091 = ~input_c[0];

  assign cgp_out[0] = 1'b0;
endmodule