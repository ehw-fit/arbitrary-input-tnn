module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050_not;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072_not;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100_not;
  wire cgp_core_101;
  wire cgp_core_103_not;
  wire cgp_core_104;
  wire cgp_core_106;
  wire cgp_core_107;

  assign cgp_core_020 = input_h[0] ^ input_i[0];
  assign cgp_core_023 = input_h[1] & input_i[1];
  assign cgp_core_027 = input_f[0] ^ cgp_core_020;
  assign cgp_core_028 = input_d[0] & cgp_core_020;
  assign cgp_core_031 = input_d[1] ^ input_c[0];
  assign cgp_core_032 = input_d[1] & cgp_core_028;
  assign cgp_core_034 = cgp_core_023 | cgp_core_032;
  assign cgp_core_035 = cgp_core_023 & cgp_core_032;
  assign cgp_core_037 = input_b[0] & input_c[0];
  assign cgp_core_039 = input_b[1] & input_c[1];
  assign cgp_core_041 = input_g[1] & cgp_core_037;
  assign cgp_core_042 = input_f[1] | input_c[1];
  assign cgp_core_044 = input_a[0] & input_g[0];
  assign cgp_core_045 = input_a[1] ^ input_b[0];
  assign cgp_core_047 = cgp_core_045 ^ input_e[1];
  assign cgp_core_048 = ~(cgp_core_045 & input_g[0]);
  assign cgp_core_050_not = ~cgp_core_042;
  assign cgp_core_052 = input_a[0] ^ input_g[0];
  assign cgp_core_053 = input_g[1] & input_g[0];
  assign cgp_core_054 = input_f[1] ^ input_h[1];
  assign cgp_core_056 = cgp_core_054 ^ input_e[1];
  assign cgp_core_057 = cgp_core_054 & cgp_core_053;
  assign cgp_core_059 = input_a[1] ^ cgp_core_052;
  assign cgp_core_060 = ~(input_e[0] & cgp_core_052);
  assign cgp_core_061 = input_e[1] ^ cgp_core_056;
  assign cgp_core_062 = ~(input_e[1] | cgp_core_056);
  assign cgp_core_063 = cgp_core_061 ^ input_d[1];
  assign cgp_core_064 = cgp_core_061 & cgp_core_060;
  assign cgp_core_065 = input_a[0] | cgp_core_064;
  assign cgp_core_066 = cgp_core_057 ^ cgp_core_065;
  assign cgp_core_067 = cgp_core_057 & cgp_core_065;
  assign cgp_core_069 = input_h[0] & input_i[0];
  assign cgp_core_071 = ~cgp_core_047;
  assign cgp_core_072_not = ~cgp_core_069;
  assign cgp_core_074 = ~input_h[1];
  assign cgp_core_076 = cgp_core_050_not & input_g[0];
  assign cgp_core_081 = input_b[1] & cgp_core_067;
  assign cgp_core_082 = cgp_core_042 ^ cgp_core_076;
  assign cgp_core_085 = ~cgp_core_081;
  assign cgp_core_086 = ~input_e[0];
  assign cgp_core_087 = ~input_d[1];
  assign cgp_core_089 = input_e[1] & cgp_core_086;
  assign cgp_core_090 = ~(cgp_core_035 ^ cgp_core_082);
  assign cgp_core_091 = cgp_core_090 & cgp_core_086;
  assign cgp_core_092 = ~cgp_core_074;
  assign cgp_core_093 = cgp_core_034 & input_c[0];
  assign cgp_core_094 = cgp_core_093 & cgp_core_091;
  assign cgp_core_095 = cgp_core_034 ^ input_h[0];
  assign cgp_core_096 = cgp_core_095 & cgp_core_091;
  assign cgp_core_097 = ~cgp_core_072_not;
  assign cgp_core_098 = ~cgp_core_031;
  assign cgp_core_099 = cgp_core_098 & cgp_core_096;
  assign cgp_core_100_not = ~cgp_core_072_not;
  assign cgp_core_101 = input_c[1] & cgp_core_096;
  assign cgp_core_103_not = ~cgp_core_027;
  assign cgp_core_104 = cgp_core_103_not & cgp_core_101;
  assign cgp_core_106 = cgp_core_027 & cgp_core_101;
  assign cgp_core_107 = input_e[0] | cgp_core_094;

  assign cgp_out[0] = 1'b0;
endmodule