module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061_not;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076_not;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017_not = ~input_d[2];
  assign cgp_core_018 = input_a[0] & input_e[0];
  assign cgp_core_022 = input_c[0] ^ input_d[1];
  assign cgp_core_023 = ~(input_e[1] & input_e[0]);
  assign cgp_core_025 = input_a[2] & input_b[2];
  assign cgp_core_027 = ~(input_a[0] ^ input_d[1]);
  assign cgp_core_031 = input_a[0] & input_a[2];
  assign cgp_core_032 = input_a[2] | input_e[1];
  assign cgp_core_033_not = ~input_c[2];
  assign cgp_core_034 = input_c[1] | input_a[2];
  assign cgp_core_035 = ~(input_d[0] & input_e[1]);
  assign cgp_core_036 = input_e[1] ^ input_c[1];
  assign cgp_core_037 = input_a[1] ^ input_c[0];
  assign cgp_core_038 = input_e[1] | input_a[1];
  assign cgp_core_039 = input_b[0] ^ input_c[1];
  assign cgp_core_040 = ~(input_d[0] ^ input_b[0]);
  assign cgp_core_041 = input_a[0] | input_b[0];
  assign cgp_core_042 = input_b[2] & input_b[2];
  assign cgp_core_043 = ~(input_e[1] ^ input_a[1]);
  assign cgp_core_044 = input_c[0] | input_c[0];
  assign cgp_core_045 = ~(input_c[0] | input_e[1]);
  assign cgp_core_046 = ~(input_a[2] & input_b[2]);
  assign cgp_core_049_not = ~input_b[1];
  assign cgp_core_050 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_051 = ~input_e[2];
  assign cgp_core_052 = input_c[0] | input_c[0];
  assign cgp_core_053 = input_a[0] ^ input_b[2];
  assign cgp_core_054 = ~(input_d[2] | input_d[2]);
  assign cgp_core_055 = ~(input_c[2] | input_d[1]);
  assign cgp_core_056 = input_e[0] | input_d[2];
  assign cgp_core_059 = cgp_core_025 & input_a[1];
  assign cgp_core_060 = ~(input_a[0] ^ input_c[0]);
  assign cgp_core_061_not = ~input_c[1];
  assign cgp_core_063 = ~(input_a[2] ^ input_d[2]);
  assign cgp_core_064 = ~(input_a[1] | input_e[0]);
  assign cgp_core_065 = ~(input_e[0] & input_d[2]);
  assign cgp_core_067 = ~(input_e[1] ^ input_a[2]);
  assign cgp_core_068 = ~(input_d[1] | input_c[2]);
  assign cgp_core_069 = input_b[2] & input_c[1];
  assign cgp_core_070 = ~(input_a[1] | input_c[1]);
  assign cgp_core_072 = input_d[0] ^ input_c[1];
  assign cgp_core_073 = input_d[0] ^ input_d[1];
  assign cgp_core_074 = input_b[0] ^ input_e[0];
  assign cgp_core_076_not = ~input_c[0];
  assign cgp_core_077 = ~(input_d[1] ^ input_e[0]);
  assign cgp_core_078 = ~(input_e[1] | input_b[2]);
  assign cgp_core_079 = ~(input_b[1] | input_b[2]);
  assign cgp_core_080 = input_b[2] & input_c[1];

  assign cgp_out[0] = cgp_core_059;
endmodule