module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018_not;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038_not;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070_not;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_076_not;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;

  assign cgp_core_018_not = ~input_f[0];
  assign cgp_core_019 = input_c[1] ^ input_g[1];
  assign cgp_core_021 = ~(input_d[0] & input_b[1]);
  assign cgp_core_022 = input_h[1] ^ input_c[1];
  assign cgp_core_023 = ~(input_e[0] | input_b[0]);
  assign cgp_core_024 = input_h[1] | input_d[1];
  assign cgp_core_026 = input_d[0] ^ input_e[1];
  assign cgp_core_028 = ~(input_h[0] & input_g[0]);
  assign cgp_core_035 = input_d[1] | input_c[0];
  assign cgp_core_037 = input_b[1] & input_c[1];
  assign cgp_core_038_not = ~input_g[0];
  assign cgp_core_042 = ~(input_d[1] & input_c[1]);
  assign cgp_core_043 = ~(input_f[0] & input_d[1]);
  assign cgp_core_045 = ~input_h[1];
  assign cgp_core_046 = ~input_b[1];
  assign cgp_core_047 = ~(input_d[0] ^ input_b[1]);
  assign cgp_core_051 = input_e[1] & input_g[1];
  assign cgp_core_052 = ~(input_a[1] | input_h[0]);
  assign cgp_core_053 = ~input_c[1];
  assign cgp_core_056 = ~(input_h[0] & input_g[1]);
  assign cgp_core_058 = input_f[1] ^ input_b[0];
  assign cgp_core_061 = ~(input_h[0] & input_f[0]);
  assign cgp_core_062 = input_c[1] | input_a[1];
  assign cgp_core_063 = input_h[0] ^ input_h[1];
  assign cgp_core_064 = cgp_core_037 | cgp_core_051;
  assign cgp_core_065 = ~input_e[1];
  assign cgp_core_066 = input_c[1] | input_g[0];
  assign cgp_core_068 = input_f[1] | cgp_core_064;
  assign cgp_core_069 = input_f[1] | cgp_core_068;
  assign cgp_core_070_not = ~input_f[1];
  assign cgp_core_072 = ~(input_h[1] ^ input_f[1]);
  assign cgp_core_074 = input_a[0] | input_d[0];
  assign cgp_core_076_not = ~cgp_core_069;
  assign cgp_core_078 = ~(input_g[1] | input_h[1]);
  assign cgp_core_079 = cgp_core_024 & input_a[1];
  assign cgp_core_080 = cgp_core_079 & cgp_core_076_not;
  assign cgp_core_081 = ~(input_a[1] | input_b[1]);
  assign cgp_core_085 = ~(input_a[1] ^ input_b[1]);
  assign cgp_core_087 = ~(input_a[0] ^ input_f[1]);
  assign cgp_core_088 = ~(input_e[0] ^ input_d[1]);
  assign cgp_core_089 = ~(input_d[1] ^ input_h[0]);
  assign cgp_core_090 = ~(input_g[0] ^ input_b[0]);
  assign cgp_core_092 = ~(input_h[1] | input_g[0]);
  assign cgp_core_093 = ~(input_d[1] ^ input_h[0]);
  assign cgp_core_094 = ~(input_e[1] & input_d[0]);
  assign cgp_core_095 = ~input_a[0];
  assign cgp_core_096 = ~(input_a[1] | input_g[1]);

  assign cgp_out[0] = cgp_core_080;
endmodule