module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053_not;
  wire cgp_core_055;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072_not;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;

  assign cgp_core_017 = input_g[0] & input_c[0];
  assign cgp_core_018 = ~input_a[1];
  assign cgp_core_019_not = ~input_b[0];
  assign cgp_core_021 = ~(cgp_core_018 ^ cgp_core_017);
  assign cgp_core_022 = ~(input_a[0] & cgp_core_021);
  assign cgp_core_024 = input_c[1] & input_g[0];
  assign cgp_core_025 = input_e[1] | input_c[0];
  assign cgp_core_026 = ~(input_e[0] & input_g[1]);
  assign cgp_core_027 = cgp_core_025 ^ cgp_core_024;
  assign cgp_core_028 = cgp_core_025 ^ input_e[1];
  assign cgp_core_029_not = ~cgp_core_028;
  assign cgp_core_030 = input_d[0] ^ input_a[0];
  assign cgp_core_032 = input_d[1] | cgp_core_027;
  assign cgp_core_034 = cgp_core_032 ^ input_f[1];
  assign cgp_core_036 = input_a[0] ^ input_d[1];
  assign cgp_core_037 = input_a[1] ^ cgp_core_036;
  assign cgp_core_038 = cgp_core_029_not | input_a[1];
  assign cgp_core_041 = ~(input_c[0] ^ cgp_core_034);
  assign cgp_core_043 = input_f[1] | input_c[0];
  assign cgp_core_045 = ~(input_e[0] ^ input_d[0]);
  assign cgp_core_046 = ~(input_b[1] | cgp_core_037);
  assign cgp_core_047 = ~(input_b[0] | input_b[0]);
  assign cgp_core_050 = ~input_c[1];
  assign cgp_core_051 = ~(cgp_core_038 & input_f[0]);
  assign cgp_core_053_not = ~input_f[0];
  assign cgp_core_055 = input_b[1] ^ input_f[1];
  assign cgp_core_061 = input_b[0] & input_a[1];
  assign cgp_core_062 = cgp_core_051 & input_g[1];
  assign cgp_core_063 = input_g[1] & input_c[0];
  assign cgp_core_065 = input_c[0] | input_b[0];
  assign cgp_core_066 = cgp_core_065 & input_f[1];
  assign cgp_core_070 = ~(input_e[1] & input_a[1]);
  assign cgp_core_071 = cgp_core_070 | input_c[1];
  assign cgp_core_072_not = ~input_b[1];
  assign cgp_core_073 = cgp_core_072_not ^ input_c[0];
  assign cgp_core_075 = input_a[1] & input_d[1];
  assign cgp_core_076 = input_b[1] & input_f[1];
  assign cgp_core_078 = input_e[0] | cgp_core_073;
  assign cgp_core_079 = ~(input_g[0] ^ cgp_core_066);
  assign cgp_core_081 = input_a[0] ^ cgp_core_078;
  assign cgp_core_082 = input_b[0] | input_a[0];

  assign cgp_out[0] = 1'b1;
endmodule