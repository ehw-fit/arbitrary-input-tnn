module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052_not;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;

  assign cgp_core_016 = ~(input_g[0] ^ input_c[1]);
  assign cgp_core_018 = input_d[1] & input_g[0];
  assign cgp_core_019 = input_c[1] & input_e[1];
  assign cgp_core_021 = ~(input_g[1] ^ input_f[0]);
  assign cgp_core_023_not = ~input_b[1];
  assign cgp_core_024 = input_e[1] & input_e[1];
  assign cgp_core_025 = input_a[1] & input_c[0];
  assign cgp_core_026 = ~(input_c[0] & input_d[1]);
  assign cgp_core_028 = input_g[1] & input_g[1];
  assign cgp_core_031 = cgp_core_019 & input_a[1];
  assign cgp_core_034 = input_d[0] | input_a[1];
  assign cgp_core_036 = ~(input_f[1] ^ input_d[0]);
  assign cgp_core_038 = ~(input_d[1] ^ input_g[0]);
  assign cgp_core_039 = input_b[1] | input_g[0];
  assign cgp_core_040 = ~(input_g[1] & input_a[1]);
  assign cgp_core_041 = ~(input_b[0] & input_a[0]);
  assign cgp_core_042 = ~(input_d[1] & input_d[0]);
  assign cgp_core_043 = ~(input_b[0] | input_f[1]);
  assign cgp_core_045 = input_g[1] ^ input_e[1];
  assign cgp_core_049 = ~input_b[1];
  assign cgp_core_050 = input_e[0] & input_b[0];
  assign cgp_core_052_not = ~input_f[1];
  assign cgp_core_054_not = ~input_d[1];
  assign cgp_core_055 = ~(input_a[1] ^ input_a[0]);
  assign cgp_core_057 = ~(input_g[1] ^ input_a[0]);
  assign cgp_core_062 = ~(input_g[0] ^ input_e[1]);
  assign cgp_core_063 = ~(input_c[1] ^ input_a[1]);
  assign cgp_core_064 = ~input_d[1];
  assign cgp_core_065 = ~input_a[1];
  assign cgp_core_068 = input_a[0] | input_f[0];
  assign cgp_core_069 = ~(input_g[0] | input_g[0]);
  assign cgp_core_070 = ~input_b[0];
  assign cgp_core_072 = input_c[0] ^ input_b[1];
  assign cgp_core_073 = ~(input_d[0] & input_b[0]);
  assign cgp_core_074 = input_c[0] ^ input_d[1];
  assign cgp_core_075 = input_e[0] & input_a[1];

  assign cgp_out[0] = cgp_core_031;
endmodule