module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_010;
  wire cgp_core_012_not;
  wire cgp_core_013;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;

  assign cgp_core_010 = ~input_d[1];
  assign cgp_core_012_not = ~input_b[1];
  assign cgp_core_013 = ~(input_a[1] | input_a[0]);
  assign cgp_core_015 = input_c[1] & input_b[0];
  assign cgp_core_016 = ~input_b[0];
  assign cgp_core_017 = ~input_d[1];
  assign cgp_core_019 = input_b[1] | input_d[1];
  assign cgp_core_020 = ~(input_c[0] | input_d[0]);
  assign cgp_core_022 = ~(input_c[0] & input_b[0]);
  assign cgp_core_025 = ~input_c[1];
  assign cgp_core_027 = input_a[0] & input_c[0];
  assign cgp_core_028_not = ~input_a[1];
  assign cgp_core_033 = ~input_a[1];
  assign cgp_core_036 = ~(input_c[0] ^ input_b[1]);
  assign cgp_core_039 = ~input_d[0];
  assign cgp_core_040 = cgp_core_033 | cgp_core_019;
  assign cgp_core_042 = input_c[1] | input_d[0];
  assign cgp_core_043 = cgp_core_040 | input_c[1];

  assign cgp_out[0] = cgp_core_043;
endmodule