module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066_not;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = ~(input_f[1] & input_c[0]);
  assign cgp_core_017 = input_c[1] & input_c[1];
  assign cgp_core_019 = input_g[0] ^ input_c[0];
  assign cgp_core_023 = input_g[0] | input_b[1];
  assign cgp_core_024 = ~(input_d[0] ^ input_c[1]);
  assign cgp_core_025 = ~input_e[0];
  assign cgp_core_026 = input_e[1] & input_g[1];
  assign cgp_core_027 = ~(input_e[1] | input_e[1]);
  assign cgp_core_030 = ~(input_d[0] & input_c[0]);
  assign cgp_core_032 = input_c[1] | input_g[1];
  assign cgp_core_036 = input_c[0] | cgp_core_032;
  assign cgp_core_038 = input_c[1] & input_g[1];
  assign cgp_core_039 = input_e[1] | cgp_core_036;
  assign cgp_core_041 = cgp_core_038 | cgp_core_026;
  assign cgp_core_042 = ~(input_g[0] | input_b[1]);
  assign cgp_core_044 = ~(input_b[0] | input_f[1]);
  assign cgp_core_045 = input_b[1] & input_f[1];
  assign cgp_core_046 = ~(input_c[0] ^ input_b[1]);
  assign cgp_core_047 = ~(input_c[1] | input_c[1]);
  assign cgp_core_049 = ~(input_c[1] ^ input_b[0]);
  assign cgp_core_050 = ~input_d[1];
  assign cgp_core_051 = ~(input_a[0] & input_e[0]);
  assign cgp_core_052 = input_f[0] | input_c[0];
  assign cgp_core_053 = input_g[0] | input_g[1];
  assign cgp_core_054 = input_a[1] & cgp_core_050;
  assign cgp_core_056 = cgp_core_045 | cgp_core_054;
  assign cgp_core_061 = ~cgp_core_056;
  assign cgp_core_062 = cgp_core_039 & cgp_core_061;
  assign cgp_core_064 = ~(input_b[1] ^ input_f[0]);
  assign cgp_core_065 = ~input_f[0];
  assign cgp_core_066_not = ~input_g[1];
  assign cgp_core_067 = input_c[0] | input_d[1];
  assign cgp_core_068 = input_e[1] & input_c[1];
  assign cgp_core_070 = ~(input_c[1] ^ input_g[0]);
  assign cgp_core_075 = input_e[1] | input_a[1];
  assign cgp_core_078 = cgp_core_062 | cgp_core_041;
  assign cgp_core_079 = cgp_core_068 | cgp_core_078;

  assign cgp_out[0] = cgp_core_079;
endmodule