module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_017_not;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036_not;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_051_not;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_077;

  assign cgp_core_015 = input_a[4] | input_a[4];
  assign cgp_core_017_not = ~input_a[6];
  assign cgp_core_019 = ~(input_a[1] | input_a[11]);
  assign cgp_core_020 = ~input_a[3];
  assign cgp_core_022 = input_a[11] | input_a[7];
  assign cgp_core_023 = input_a[9] | input_a[6];
  assign cgp_core_024 = input_a[6] & input_a[8];
  assign cgp_core_026 = input_a[4] & input_a[1];
  assign cgp_core_028 = ~(input_a[1] ^ input_a[3]);
  assign cgp_core_029_not = ~input_a[9];
  assign cgp_core_031 = ~(input_a[2] & input_a[8]);
  assign cgp_core_032 = ~(input_a[4] & input_a[10]);
  assign cgp_core_033 = ~input_a[3];
  assign cgp_core_036_not = ~input_a[4];
  assign cgp_core_037 = ~(input_a[2] | input_a[5]);
  assign cgp_core_040 = input_a[10] | input_a[0];
  assign cgp_core_045 = ~(input_a[11] & input_a[9]);
  assign cgp_core_046 = ~(input_a[10] ^ input_a[1]);
  assign cgp_core_047 = ~input_a[6];
  assign cgp_core_049 = input_a[5] | input_a[11];
  assign cgp_core_051_not = ~input_a[9];
  assign cgp_core_054 = input_a[5] | input_a[8];
  assign cgp_core_055 = input_a[8] ^ input_a[0];
  assign cgp_core_057 = input_a[8] | input_a[2];
  assign cgp_core_058 = input_a[1] ^ input_a[10];
  assign cgp_core_060 = input_a[7] & input_a[1];
  assign cgp_core_062 = input_a[4] & input_a[6];
  assign cgp_core_063 = ~(input_a[9] & input_a[0]);
  assign cgp_core_064 = ~(input_a[3] ^ input_a[10]);
  assign cgp_core_066 = ~input_a[0];
  assign cgp_core_070 = ~(input_a[3] & input_a[1]);
  assign cgp_core_071 = ~input_a[2];
  assign cgp_core_073 = input_a[8] ^ input_a[6];
  assign cgp_core_077 = ~(input_a[4] | input_a[11]);

  assign cgp_out[0] = input_a[7];
  assign cgp_out[1] = input_a[1];
  assign cgp_out[2] = cgp_core_047;
  assign cgp_out[3] = input_a[6];
endmodule