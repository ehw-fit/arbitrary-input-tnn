module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_022_not;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047_not;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060_not;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068_not;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = input_d[1] | input_b[1];
  assign cgp_core_018 = input_a[0] | input_f[1];
  assign cgp_core_021 = input_f[0] | input_f[0];
  assign cgp_core_022_not = ~input_d[0];
  assign cgp_core_026 = ~(input_b[1] ^ input_f[0]);
  assign cgp_core_029 = ~input_f[1];
  assign cgp_core_030 = ~(input_f[0] ^ input_g[1]);
  assign cgp_core_031 = ~(input_g[1] | input_b[1]);
  assign cgp_core_034 = input_e[0] & input_d[0];
  assign cgp_core_035 = input_f[1] | input_a[1];
  assign cgp_core_036 = input_f[0] | input_b[1];
  assign cgp_core_038 = ~(input_f[1] | input_a[1]);
  assign cgp_core_039 = ~(input_c[1] | input_c[1]);
  assign cgp_core_042 = input_d[0] ^ input_b[1];
  assign cgp_core_043 = input_e[1] & input_d[1];
  assign cgp_core_044 = ~(input_d[1] & input_d[0]);
  assign cgp_core_045 = ~input_d[1];
  assign cgp_core_047_not = ~input_f[0];
  assign cgp_core_048 = input_a[0] & input_a[0];
  assign cgp_core_049 = input_d[1] & input_c[1];
  assign cgp_core_050 = input_a[1] ^ input_g[0];
  assign cgp_core_051 = input_e[0] & input_g[1];
  assign cgp_core_052 = input_c[0] | input_f[1];
  assign cgp_core_054 = ~(input_b[1] | input_d[1]);
  assign cgp_core_055 = input_b[1] ^ input_b[1];
  assign cgp_core_056 = ~(input_g[1] & input_e[1]);
  assign cgp_core_057 = input_f[1] | input_b[1];
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = input_a[1] & cgp_core_058;
  assign cgp_core_060_not = ~input_c[1];
  assign cgp_core_061 = input_d[1] | input_f[1];
  assign cgp_core_063 = input_a[0] & input_g[0];
  assign cgp_core_065 = ~input_b[0];
  assign cgp_core_066 = ~input_f[1];
  assign cgp_core_067 = ~(input_b[1] & input_f[1]);
  assign cgp_core_068_not = ~input_a[0];
  assign cgp_core_069 = ~(input_a[1] & input_f[0]);
  assign cgp_core_071 = input_c[1] ^ input_d[0];
  assign cgp_core_074 = ~(input_e[0] ^ input_e[1]);
  assign cgp_core_075 = input_d[0] | input_c[1];
  assign cgp_core_078 = input_f[1] ^ input_b[0];
  assign cgp_core_079 = ~(input_g[0] ^ input_f[0]);

  assign cgp_out[0] = cgp_core_059;
endmodule