module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_056_not;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061_not;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087_not;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;

  assign cgp_core_016 = input_a[1] | input_a[2];
  assign cgp_core_017 = input_a[1] & input_a[2];
  assign cgp_core_019 = input_a[0] & cgp_core_016;
  assign cgp_core_020 = cgp_core_017 | cgp_core_019;
  assign cgp_core_022 = ~(input_a[3] & input_a[4]);
  assign cgp_core_023 = input_a[3] & input_a[4];
  assign cgp_core_024 = ~(input_a[5] & input_a[6]);
  assign cgp_core_025 = input_a[5] & input_a[6];
  assign cgp_core_026 = cgp_core_022 ^ cgp_core_024;
  assign cgp_core_027 = ~input_a[2];
  assign cgp_core_028 = ~(cgp_core_023 & cgp_core_025);
  assign cgp_core_035 = ~(cgp_core_020 & cgp_core_028);
  assign cgp_core_037 = cgp_core_035 ^ cgp_core_026;
  assign cgp_core_038 = input_a[5] & input_a[6];
  assign cgp_core_039 = cgp_core_020 | cgp_core_038;
  assign cgp_core_042 = cgp_core_023 | cgp_core_039;
  assign cgp_core_043 = input_a[8] ^ input_a[3];
  assign cgp_core_044 = ~(input_a[7] & input_a[12]);
  assign cgp_core_045 = input_a[8] ^ input_a[9];
  assign cgp_core_046 = input_a[8] & input_a[9];
  assign cgp_core_047 = input_a[7] ^ cgp_core_045;
  assign cgp_core_048 = input_a[7] & cgp_core_045;
  assign cgp_core_049 = cgp_core_046 | cgp_core_048;
  assign cgp_core_051 = input_a[11] ^ input_a[12];
  assign cgp_core_052 = ~(input_a[12] & input_a[5]);
  assign cgp_core_054 = ~(input_a[13] & input_a[10]);
  assign cgp_core_056_not = ~input_a[0];
  assign cgp_core_058 = input_a[1] & input_a[13];
  assign cgp_core_059 = input_a[11] & input_a[12];
  assign cgp_core_060 = ~input_a[3];
  assign cgp_core_061_not = ~input_a[0];
  assign cgp_core_062 = cgp_core_047 ^ input_a[10];
  assign cgp_core_063 = cgp_core_047 & input_a[10];
  assign cgp_core_064 = cgp_core_049 ^ cgp_core_059;
  assign cgp_core_065 = cgp_core_049 & cgp_core_059;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_070 = ~(input_a[0] | input_a[13]);
  assign cgp_core_074 = ~(input_a[8] ^ input_a[13]);
  assign cgp_core_075 = input_a[13] & cgp_core_062;
  assign cgp_core_076 = cgp_core_037 ^ cgp_core_066;
  assign cgp_core_077 = cgp_core_037 & cgp_core_066;
  assign cgp_core_078 = cgp_core_076 ^ cgp_core_075;
  assign cgp_core_079 = cgp_core_076 & cgp_core_075;
  assign cgp_core_080 = cgp_core_077 | cgp_core_079;
  assign cgp_core_081 = cgp_core_042 ^ cgp_core_068;
  assign cgp_core_082 = cgp_core_042 & cgp_core_068;
  assign cgp_core_083 = cgp_core_081 ^ cgp_core_080;
  assign cgp_core_084 = cgp_core_081 & cgp_core_080;
  assign cgp_core_085 = cgp_core_082 | cgp_core_084;
  assign cgp_core_087_not = ~input_a[1];
  assign cgp_core_088 = input_a[5] & input_a[12];
  assign cgp_core_089 = input_a[2] | input_a[10];
  assign cgp_core_090 = input_a[9] & input_a[1];

  assign cgp_out[0] = cgp_core_051;
  assign cgp_out[1] = cgp_core_078;
  assign cgp_out[2] = cgp_core_083;
  assign cgp_out[3] = cgp_core_085;
endmodule