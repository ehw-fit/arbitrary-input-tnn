module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018_not;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;

  assign cgp_core_011 = ~input_b[0];
  assign cgp_core_014 = input_a[1] & input_b[1];
  assign cgp_core_015 = ~input_b[2];
  assign cgp_core_017 = cgp_core_014 | input_a[2];
  assign cgp_core_018_not = ~input_b[2];
  assign cgp_core_019 = ~input_a[1];
  assign cgp_core_020 = input_b[0] | input_a[2];
  assign cgp_core_022 = input_b[2] | cgp_core_017;
  assign cgp_core_024 = ~input_a[1];
  assign cgp_core_029 = ~input_c[2];
  assign cgp_core_030 = ~(input_a[2] | input_c[1]);
  assign cgp_core_032 = input_c[0] ^ input_a[0];
  assign cgp_core_033 = input_c[0] | input_b[2];
  assign cgp_core_034 = input_c[2] | input_a[0];
  assign cgp_core_035 = input_a[0] ^ input_a[0];
  assign cgp_core_037 = input_b[0] ^ input_a[1];
  assign cgp_core_038 = ~input_b[1];
  assign cgp_core_039 = input_b[1] & input_a[1];

  assign cgp_out[0] = cgp_core_022;
endmodule