module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_081;
  wire cgp_core_082_not;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;
  wire cgp_core_097;
  wire cgp_core_100;
  wire cgp_core_103;
  wire cgp_core_109_not;
  wire cgp_core_110;

  assign cgp_core_021 = input_h[0] & input_i[0];
  assign cgp_core_022 = input_h[1] ^ input_i[1];
  assign cgp_core_023 = input_i[1] & input_c[1];
  assign cgp_core_026 = cgp_core_023 | input_g[1];
  assign cgp_core_029 = input_d[1] ^ input_a[1];
  assign cgp_core_030 = ~(input_d[1] ^ input_f[1]);
  assign cgp_core_031 = ~(input_a[1] ^ input_d[0]);
  assign cgp_core_032 = input_i[1] & input_f[0];
  assign cgp_core_033 = input_d[1] | input_e[0];
  assign cgp_core_035 = ~(cgp_core_026 & input_a[1]);
  assign cgp_core_036_not = ~input_c[0];
  assign cgp_core_038 = input_c[0] ^ input_c[1];
  assign cgp_core_039 = input_d[0] | input_d[1];
  assign cgp_core_043 = ~(input_a[0] | input_d[0]);
  assign cgp_core_044 = input_a[0] & input_c[1];
  assign cgp_core_045 = input_a[1] ^ input_b[0];
  assign cgp_core_046 = input_a[1] & cgp_core_038;
  assign cgp_core_047 = ~(cgp_core_045 ^ input_d[1]);
  assign cgp_core_048 = input_f[1] & cgp_core_044;
  assign cgp_core_049 = ~(cgp_core_046 | input_i[1]);
  assign cgp_core_052 = input_f[0] & input_g[0];
  assign cgp_core_053 = input_f[0] | input_g[0];
  assign cgp_core_056 = ~input_b[0];
  assign cgp_core_058 = ~(input_a[0] & input_h[0]);
  assign cgp_core_059 = input_b[1] & cgp_core_052;
  assign cgp_core_060 = input_e[0] & cgp_core_052;
  assign cgp_core_061 = input_e[1] | input_f[1];
  assign cgp_core_062 = input_g[1] & cgp_core_056;
  assign cgp_core_063 = input_a[1] ^ cgp_core_060;
  assign cgp_core_064 = input_d[1] & input_i[0];
  assign cgp_core_065 = ~(cgp_core_062 ^ cgp_core_064);
  assign cgp_core_066 = ~input_c[0];
  assign cgp_core_067 = input_a[0] & cgp_core_065;
  assign cgp_core_068 = cgp_core_043 ^ cgp_core_059;
  assign cgp_core_069 = cgp_core_043 ^ cgp_core_059;
  assign cgp_core_070 = ~(input_i[1] | cgp_core_063);
  assign cgp_core_071 = cgp_core_047 & input_g[0];
  assign cgp_core_072 = ~(cgp_core_070 ^ cgp_core_069);
  assign cgp_core_073 = input_g[1] & cgp_core_069;
  assign cgp_core_074 = input_g[1] | cgp_core_073;
  assign cgp_core_076 = input_f[1] & cgp_core_066;
  assign cgp_core_081 = input_b[1] & input_h[0];
  assign cgp_core_082_not = ~cgp_core_067;
  assign cgp_core_085 = ~input_f[0];
  assign cgp_core_087 = ~input_h[0];
  assign cgp_core_088 = cgp_core_035 & input_a[1];
  assign cgp_core_089 = input_d[1] | input_h[0];
  assign cgp_core_090 = ~(cgp_core_035 ^ cgp_core_082_not);
  assign cgp_core_091 = ~input_e[1];
  assign cgp_core_093 = input_g[1] & input_i[1];
  assign cgp_core_097 = ~cgp_core_072;
  assign cgp_core_100 = ~(input_a[0] ^ input_a[1]);
  assign cgp_core_103 = input_d[0] & input_h[0];
  assign cgp_core_109_not = ~input_c[0];
  assign cgp_core_110 = input_g[1] | cgp_core_109_not;

  assign cgp_out[0] = 1'b0;
endmodule