module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_010;
  wire cgp_core_013_not;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_026;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_043;

  assign cgp_core_010 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_013_not = ~input_a[0];
  assign cgp_core_014 = ~(input_b[1] | input_d[0]);
  assign cgp_core_015 = input_d[0] & input_a[1];
  assign cgp_core_016 = input_a[1] | input_a[1];
  assign cgp_core_017 = input_d[0] | input_b[0];
  assign cgp_core_020 = ~(input_b[1] ^ input_b[0]);
  assign cgp_core_021 = input_c[0] | input_b[1];
  assign cgp_core_022 = input_d[1] | input_c[0];
  assign cgp_core_023 = ~input_a[1];
  assign cgp_core_024_not = ~input_d[0];
  assign cgp_core_026 = input_d[0] ^ input_d[1];
  assign cgp_core_031 = ~input_b[0];
  assign cgp_core_032 = ~input_c[1];
  assign cgp_core_034 = ~(input_a[0] | input_d[1]);
  assign cgp_core_035 = ~input_a[0];
  assign cgp_core_039 = ~(input_b[0] & input_d[0]);
  assign cgp_core_040 = input_c[1] | input_d[1];
  assign cgp_core_041_not = ~input_d[1];
  assign cgp_core_042 = input_b[0] | input_b[1];
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;

  assign cgp_out[0] = cgp_core_043;
endmodule