module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_014 = input_e[1] & input_d[0];
  assign cgp_core_015 = input_e[0] & input_d[0];
  assign cgp_core_016 = input_a[0] | input_d[0];
  assign cgp_core_017 = ~input_b[1];
  assign cgp_core_018 = input_a[1] | cgp_core_015;
  assign cgp_core_019 = ~(input_e[1] & input_d[1]);
  assign cgp_core_020 = input_f[1] & input_c[0];
  assign cgp_core_021 = input_c[1] ^ input_f[0];
  assign cgp_core_023 = input_f[1] & input_d[1];
  assign cgp_core_024 = ~input_c[1];
  assign cgp_core_025 = ~(input_c[0] | input_c[1]);
  assign cgp_core_029 = ~(input_a[1] ^ input_e[0]);
  assign cgp_core_030 = ~input_e[1];
  assign cgp_core_031 = ~input_b[1];
  assign cgp_core_032 = ~input_c[1];
  assign cgp_core_033 = ~input_e[1];
  assign cgp_core_035 = input_f[1] & input_f[0];
  assign cgp_core_036 = input_d[1] | input_c[1];
  assign cgp_core_037 = input_c[1] & input_a[1];
  assign cgp_core_038 = input_f[1] ^ input_c[1];
  assign cgp_core_039 = input_f[0] ^ input_e[0];
  assign cgp_core_041 = ~(input_c[1] ^ input_c[0]);
  assign cgp_core_045 = ~(input_b[0] & input_f[1]);
  assign cgp_core_046 = input_d[1] | cgp_core_018;
  assign cgp_core_048 = ~input_c[1];
  assign cgp_core_049 = ~(input_e[1] ^ input_d[1]);
  assign cgp_core_050 = input_b[0] & input_d[1];
  assign cgp_core_053 = ~(input_d[0] ^ input_a[1]);
  assign cgp_core_054 = ~(input_c[0] & input_c[0]);
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_061 = input_b[1] ^ input_d[0];
  assign cgp_core_063 = ~(input_d[1] | input_e[1]);
  assign cgp_core_066 = ~(input_b[0] | input_a[0]);
  assign cgp_core_067 = input_a[0] & input_c[0];
  assign cgp_core_068 = cgp_core_058 | cgp_core_046;
  assign cgp_core_069 = input_e[1] | cgp_core_068;
  assign cgp_core_070 = input_c[1] | cgp_core_067;
  assign cgp_core_071 = input_f[1] | cgp_core_070;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;

  assign cgp_out[0] = cgp_core_072;
endmodule