module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021_not;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_026_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;

  assign cgp_core_017 = ~(input_a[1] ^ input_c[0]);
  assign cgp_core_018 = ~input_d[0];
  assign cgp_core_020 = input_c[0] ^ input_b[1];
  assign cgp_core_021_not = ~input_d[0];
  assign cgp_core_022 = input_e[1] ^ input_c[1];
  assign cgp_core_023 = input_c[2] & input_e[2];
  assign cgp_core_026_not = ~input_e[0];
  assign cgp_core_028 = ~input_d[1];
  assign cgp_core_029 = ~(input_c[0] & input_e[1]);
  assign cgp_core_030 = input_a[1] | input_c[1];
  assign cgp_core_031 = input_e[0] ^ input_d[0];
  assign cgp_core_032 = ~input_d[0];
  assign cgp_core_033 = ~(input_d[1] ^ input_e[2]);
  assign cgp_core_035 = input_b[0] & input_a[2];
  assign cgp_core_036 = input_d[2] | input_b[2];
  assign cgp_core_037 = input_b[1] & input_d[0];
  assign cgp_core_041 = ~(input_e[2] ^ input_c[2]);
  assign cgp_core_042 = ~(input_d[2] & input_a[2]);
  assign cgp_core_044 = input_c[1] & input_e[0];
  assign cgp_core_045_not = ~input_e[2];
  assign cgp_core_046 = ~(input_c[1] | input_b[1]);
  assign cgp_core_047 = ~(input_b[2] ^ input_d[0]);
  assign cgp_core_049 = input_c[0] & input_d[2];
  assign cgp_core_052 = ~(input_d[0] & input_c[2]);
  assign cgp_core_053 = ~(input_b[1] ^ input_c[0]);
  assign cgp_core_055 = ~(input_c[1] & input_a[0]);
  assign cgp_core_057 = input_b[0] ^ input_a[2];
  assign cgp_core_058 = input_e[2] ^ input_c[2];
  assign cgp_core_059 = input_b[2] ^ input_c[1];
  assign cgp_core_060 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_063 = input_a[0] ^ input_c[1];
  assign cgp_core_064 = ~(input_b[2] | input_d[0]);
  assign cgp_core_067 = input_e[1] & input_a[1];
  assign cgp_core_068 = input_b[2] & input_c[2];
  assign cgp_core_069 = ~(input_d[2] | input_c[0]);
  assign cgp_core_070 = ~input_d[2];
  assign cgp_core_071 = input_e[0] & input_e[1];
  assign cgp_core_072 = ~(input_e[2] | input_d[2]);
  assign cgp_core_073 = ~(input_c[2] ^ input_d[2]);
  assign cgp_core_074_not = ~input_a[1];
  assign cgp_core_075 = input_a[2] ^ input_d[1];
  assign cgp_core_076 = ~(input_c[2] & input_e[0]);
  assign cgp_core_077 = input_a[0] ^ input_d[0];

  assign cgp_out[0] = cgp_core_042;
endmodule