module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_056_not;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_080;
  wire cgp_core_082_not;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_099;
  wire cgp_core_101;
  wire cgp_core_103;
  wire cgp_core_104;

  assign cgp_core_020 = input_h[0] ^ input_i[0];
  assign cgp_core_021 = input_b[1] | input_i[0];
  assign cgp_core_022 = input_h[1] ^ input_i[1];
  assign cgp_core_024 = input_h[0] ^ cgp_core_021;
  assign cgp_core_028 = ~(input_d[0] ^ input_h[1]);
  assign cgp_core_029 = input_d[1] ^ cgp_core_024;
  assign cgp_core_030 = input_d[1] & cgp_core_024;
  assign cgp_core_032 = cgp_core_029 & cgp_core_028;
  assign cgp_core_033 = input_c[1] | input_d[1];
  assign cgp_core_034_not = ~cgp_core_033;
  assign cgp_core_037 = input_b[0] & input_c[0];
  assign cgp_core_038 = input_b[1] ^ input_c[1];
  assign cgp_core_040 = input_g[0] ^ input_h[1];
  assign cgp_core_041 = cgp_core_038 & input_i[0];
  assign cgp_core_043 = input_a[0] ^ input_d[0];
  assign cgp_core_045 = input_e[1] ^ cgp_core_040;
  assign cgp_core_046 = ~input_a[1];
  assign cgp_core_047 = input_i[1] ^ input_h[1];
  assign cgp_core_049 = ~(cgp_core_046 | cgp_core_045);
  assign cgp_core_052 = ~(input_f[1] & input_g[0]);
  assign cgp_core_053 = input_f[0] & input_f[1];
  assign cgp_core_056_not = ~cgp_core_053;
  assign cgp_core_060 = input_e[0] & cgp_core_052;
  assign cgp_core_061 = input_e[1] ^ cgp_core_056_not;
  assign cgp_core_062 = ~input_e[1];
  assign cgp_core_063 = cgp_core_061 ^ input_b[0];
  assign cgp_core_064 = input_b[1] & cgp_core_060;
  assign cgp_core_071 = cgp_core_047 & cgp_core_063;
  assign cgp_core_074 = input_g[0] ^ input_i[0];
  assign cgp_core_080 = input_a[0] ^ input_f[1];
  assign cgp_core_082_not = ~input_g[1];
  assign cgp_core_083 = cgp_core_080 & input_g[0];
  assign cgp_core_084 = input_d[0] & input_f[1];
  assign cgp_core_085 = ~cgp_core_084;
  assign cgp_core_087 = ~cgp_core_082_not;
  assign cgp_core_092 = ~input_b[1];
  assign cgp_core_093 = cgp_core_034_not & cgp_core_092;
  assign cgp_core_094 = ~(input_c[0] & input_c[1]);
  assign cgp_core_096 = input_c[1] & input_e[1];
  assign cgp_core_097 = ~input_c[1];
  assign cgp_core_099 = ~(input_c[0] & cgp_core_096);
  assign cgp_core_101 = input_i[0] & cgp_core_096;
  assign cgp_core_103 = ~input_b[1];
  assign cgp_core_104 = cgp_core_103 & cgp_core_101;

  assign cgp_out[0] = 1'b0;
endmodule