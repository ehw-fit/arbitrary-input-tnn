module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_015;
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_012 = input_a[1] | input_d[1];
  assign cgp_core_013 = ~(input_e[0] | input_d[0]);
  assign cgp_core_015 = ~input_a[1];
  assign cgp_core_018 = input_d[1] | input_b[1];
  assign cgp_core_019_not = ~input_b[1];
  assign cgp_core_021 = input_b[1] ^ input_e[0];
  assign cgp_core_022 = input_c[1] & input_e[1];
  assign cgp_core_024 = input_a[1] & input_a[0];
  assign cgp_core_025 = cgp_core_022 | cgp_core_024;
  assign cgp_core_026 = ~(input_e[0] ^ input_e[1]);
  assign cgp_core_027_not = ~input_b[0];
  assign cgp_core_028 = input_e[0] ^ input_e[0];
  assign cgp_core_029 = input_a[1] & input_c[0];
  assign cgp_core_033 = cgp_core_025 | cgp_core_029;
  assign cgp_core_035 = ~(input_a[0] | input_a[0]);
  assign cgp_core_036 = ~(input_d[1] & input_d[0]);
  assign cgp_core_037 = ~cgp_core_033;
  assign cgp_core_038 = cgp_core_018 & cgp_core_037;
  assign cgp_core_039 = ~(input_e[0] | input_a[0]);
  assign cgp_core_040 = ~(input_a[0] ^ input_e[1]);
  assign cgp_core_042 = input_e[0] ^ input_b[0];
  assign cgp_core_045 = input_c[0] ^ input_d[1];
  assign cgp_core_046 = input_d[0] & input_b[1];
  assign cgp_core_047_not = ~input_e[0];
  assign cgp_core_049 = ~input_c[1];
  assign cgp_core_050 = ~input_b[0];
  assign cgp_core_051 = ~(input_c[1] & input_c[1]);
  assign cgp_core_053 = input_c[0] | input_b[0];
  assign cgp_core_054 = ~input_a[1];

  assign cgp_out[0] = cgp_core_038;
endmodule