module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027_not;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052_not;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090_not;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_101;
  wire cgp_core_102;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_110;

  assign cgp_core_022 = input_h[1] ^ input_i[1];
  assign cgp_core_023 = input_h[1] & input_i[1];
  assign cgp_core_025 = input_h[0] ^ input_a[1];
  assign cgp_core_027_not = ~input_f[1];
  assign cgp_core_028_not = ~input_c[1];
  assign cgp_core_029 = input_d[1] ^ cgp_core_022;
  assign cgp_core_030 = input_d[1] & cgp_core_022;
  assign cgp_core_032 = input_a[0] | input_i[1];
  assign cgp_core_034 = cgp_core_023 | cgp_core_030;
  assign cgp_core_037 = input_i[1] & input_e[1];
  assign cgp_core_038 = input_b[1] | input_c[1];
  assign cgp_core_039 = ~(input_i[0] & input_d[1]);
  assign cgp_core_040 = cgp_core_038 ^ input_b[0];
  assign cgp_core_041 = cgp_core_038 & input_b[0];
  assign cgp_core_045 = input_a[1] ^ cgp_core_040;
  assign cgp_core_046 = input_a[1] & cgp_core_040;
  assign cgp_core_047 = cgp_core_045 ^ input_g[0];
  assign cgp_core_048 = cgp_core_045 & input_g[0];
  assign cgp_core_049 = cgp_core_046 | cgp_core_048;
  assign cgp_core_050 = cgp_core_041 | cgp_core_049;
  assign cgp_core_051 = cgp_core_041 & cgp_core_049;
  assign cgp_core_052_not = ~input_c[0];
  assign cgp_core_053 = ~input_c[0];
  assign cgp_core_054 = input_f[1] | input_g[1];
  assign cgp_core_055 = input_f[1] & input_g[1];
  assign cgp_core_057 = input_d[1] | input_g[0];
  assign cgp_core_059 = ~(input_g[0] ^ input_d[1]);
  assign cgp_core_060 = input_d[0] | input_b[0];
  assign cgp_core_061 = input_e[1] | cgp_core_054;
  assign cgp_core_062 = input_e[1] & cgp_core_054;
  assign cgp_core_064 = ~input_h[0];
  assign cgp_core_066 = cgp_core_055 | cgp_core_062;
  assign cgp_core_067 = input_b[1] & input_c[1];
  assign cgp_core_068 = ~(input_h[0] | input_i[0]);
  assign cgp_core_069 = input_c[0] & input_e[0];
  assign cgp_core_070 = cgp_core_047 | cgp_core_061;
  assign cgp_core_071 = cgp_core_047 & cgp_core_061;
  assign cgp_core_073 = cgp_core_070 & cgp_core_069;
  assign cgp_core_074 = cgp_core_071 | cgp_core_073;
  assign cgp_core_075 = cgp_core_050 | cgp_core_066;
  assign cgp_core_077 = cgp_core_075 | cgp_core_074;
  assign cgp_core_078 = cgp_core_075 & cgp_core_074;
  assign cgp_core_079 = cgp_core_066 | cgp_core_078;
  assign cgp_core_080 = cgp_core_051 | cgp_core_067;
  assign cgp_core_082 = cgp_core_080 | cgp_core_079;
  assign cgp_core_083 = input_a[0] & input_f[0];
  assign cgp_core_085 = ~(input_b[0] & input_d[0]);
  assign cgp_core_086 = input_f[1] & input_f[1];
  assign cgp_core_087 = ~(input_a[0] | input_d[1]);
  assign cgp_core_089 = input_g[1] | input_e[0];
  assign cgp_core_090_not = ~cgp_core_082;
  assign cgp_core_092 = ~cgp_core_077;
  assign cgp_core_093 = cgp_core_034 & cgp_core_092;
  assign cgp_core_095 = ~(cgp_core_034 ^ cgp_core_077);
  assign cgp_core_096 = cgp_core_095 & cgp_core_090_not;
  assign cgp_core_097 = ~(input_h[1] & input_d[1]);
  assign cgp_core_099 = cgp_core_029 & cgp_core_096;
  assign cgp_core_100 = ~(input_a[0] | input_a[1]);
  assign cgp_core_101 = cgp_core_100 & cgp_core_096;
  assign cgp_core_102 = input_g[1] ^ input_e[1];
  assign cgp_core_105 = input_d[0] & input_b[1];
  assign cgp_core_106 = input_i[0] & cgp_core_101;
  assign cgp_core_107 = cgp_core_099 | cgp_core_093;
  assign cgp_core_110 = cgp_core_107 | cgp_core_106;

  assign cgp_out[0] = cgp_core_110;
endmodule