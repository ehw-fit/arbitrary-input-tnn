module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_081_not;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_088;
  wire cgp_core_095_not;

  assign cgp_core_019 = ~input_e[1];
  assign cgp_core_020 = ~(input_f[0] | input_c[0]);
  assign cgp_core_022 = ~(cgp_core_020 & input_h[0]);
  assign cgp_core_023 = ~input_d[1];
  assign cgp_core_024 = input_c[0] | input_g[1];
  assign cgp_core_025_not = ~input_d[0];
  assign cgp_core_026 = input_a[0] ^ input_e[0];
  assign cgp_core_027 = ~input_d[0];
  assign cgp_core_028 = input_a[1] & input_e[0];
  assign cgp_core_029 = input_b[1] ^ cgp_core_026;
  assign cgp_core_031 = ~(cgp_core_028 | input_h[1]);
  assign cgp_core_032 = ~(input_d[1] | input_a[1]);
  assign cgp_core_035 = input_a[1] & input_f[0];
  assign cgp_core_036 = input_d[1] & input_d[0];
  assign cgp_core_037 = ~(input_a[1] ^ input_h[1]);
  assign cgp_core_039 = input_g[1] & input_f[0];
  assign cgp_core_040 = cgp_core_037 | input_a[0];
  assign cgp_core_041 = input_e[0] ^ input_g[0];
  assign cgp_core_042 = input_h[1] | input_c[1];
  assign cgp_core_043 = ~(input_c[0] | input_h[1]);
  assign cgp_core_045 = cgp_core_043 & input_b[0];
  assign cgp_core_046 = cgp_core_043 | input_f[0];
  assign cgp_core_050 = ~cgp_core_025_not;
  assign cgp_core_052 = ~(input_b[0] | input_g[1]);
  assign cgp_core_054 = input_h[0] | input_b[1];
  assign cgp_core_055 = ~input_c[1];
  assign cgp_core_056 = input_h[0] | input_e[1];
  assign cgp_core_058 = ~(input_b[0] & input_c[1]);
  assign cgp_core_060 = ~input_g[1];
  assign cgp_core_061 = ~(cgp_core_058 ^ input_c[0]);
  assign cgp_core_062 = input_h[0] & input_c[1];
  assign cgp_core_065 = ~input_d[1];
  assign cgp_core_067 = input_g[0] ^ input_f[0];
  assign cgp_core_068 = input_b[0] & input_h[0];
  assign cgp_core_069 = input_h[0] ^ input_a[0];
  assign cgp_core_071 = input_g[1] ^ input_e[0];
  assign cgp_core_072 = input_h[0] & input_b[0];
  assign cgp_core_073 = ~input_h[1];
  assign cgp_core_074_not = ~input_e[0];
  assign cgp_core_075 = input_b[0] & input_b[1];
  assign cgp_core_076 = ~input_e[0];
  assign cgp_core_077 = ~(input_b[0] | input_b[1]);
  assign cgp_core_079 = cgp_core_056 & input_e[0];
  assign cgp_core_081_not = ~cgp_core_056;
  assign cgp_core_082 = input_e[1] & input_e[1];
  assign cgp_core_083 = ~(input_d[1] | input_b[0]);
  assign cgp_core_084 = ~(input_g[0] ^ input_d[1]);
  assign cgp_core_085 = cgp_core_084 | input_b[0];
  assign cgp_core_088 = input_a[0] ^ input_b[1];
  assign cgp_core_095_not = ~input_f[0];

  assign cgp_out[0] = 1'b1;
endmodule