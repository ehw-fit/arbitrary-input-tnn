module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_080_not;

  assign cgp_core_017 = input_c[0] ^ input_c[1];
  assign cgp_core_018 = input_a[0] & input_c[0];
  assign cgp_core_019 = input_b[1] | input_c[1];
  assign cgp_core_020 = input_b[1] & input_c[1];
  assign cgp_core_021 = cgp_core_019 | cgp_core_018;
  assign cgp_core_022 = cgp_core_019 & cgp_core_018;
  assign cgp_core_023 = cgp_core_020 | cgp_core_022;
  assign cgp_core_024 = input_b[2] | input_c[2];
  assign cgp_core_025 = input_b[2] & input_c[2];
  assign cgp_core_026 = cgp_core_024 | cgp_core_023;
  assign cgp_core_027 = cgp_core_024 & cgp_core_023;
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_029 = input_b[0] | input_b[2];
  assign cgp_core_031 = input_d[1] | input_e[1];
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_036 = input_d[2] | input_e[2];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038 = cgp_core_036 | cgp_core_032;
  assign cgp_core_039 = cgp_core_036 & input_e[1];
  assign cgp_core_040 = cgp_core_037 | cgp_core_039;
  assign cgp_core_041 = input_e[0] | input_c[0];
  assign cgp_core_042 = ~(input_c[2] & input_d[0]);
  assign cgp_core_043 = ~input_a[0];
  assign cgp_core_044 = cgp_core_021 & cgp_core_031;
  assign cgp_core_045 = input_c[0] & input_e[0];
  assign cgp_core_046 = ~input_c[1];
  assign cgp_core_048 = cgp_core_026 | cgp_core_038;
  assign cgp_core_049 = cgp_core_026 & cgp_core_038;
  assign cgp_core_050 = cgp_core_048 | cgp_core_044;
  assign cgp_core_051 = cgp_core_048 & cgp_core_044;
  assign cgp_core_052 = cgp_core_049 | cgp_core_051;
  assign cgp_core_053 = cgp_core_028 | cgp_core_040;
  assign cgp_core_054 = ~(input_a[0] ^ input_b[1]);
  assign cgp_core_055 = cgp_core_053 | cgp_core_052;
  assign cgp_core_056 = ~(input_c[0] | input_e[0]);
  assign cgp_core_058 = input_b[1] ^ input_b[0];
  assign cgp_core_059 = input_e[0] ^ input_d[1];
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_063 = ~cgp_core_050;
  assign cgp_core_064 = input_a[2] & cgp_core_063;
  assign cgp_core_066 = ~(input_a[2] ^ cgp_core_050);
  assign cgp_core_067 = cgp_core_066 & cgp_core_061;
  assign cgp_core_068 = ~input_a[0];
  assign cgp_core_069_not = ~input_e[2];
  assign cgp_core_072 = input_a[0] & cgp_core_067;
  assign cgp_core_075 = input_a[1] & cgp_core_072;
  assign cgp_core_076 = ~(input_e[1] | input_a[2]);
  assign cgp_core_077 = input_a[0] | input_e[1];
  assign cgp_core_079 = cgp_core_075 | cgp_core_064;
  assign cgp_core_080_not = ~input_a[1];

  assign cgp_out[0] = cgp_core_079;
endmodule