module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_080;

  assign cgp_core_020 = input_a[1] & input_b[1];
  assign cgp_core_024 = input_a[2] ^ input_b[2];
  assign cgp_core_025 = input_a[2] & input_b[2];
  assign cgp_core_026 = cgp_core_024 ^ cgp_core_020;
  assign cgp_core_027 = cgp_core_024 & cgp_core_020;
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_029 = ~(input_a[0] ^ input_a[2]);
  assign cgp_core_030 = input_a[1] ^ input_b[2];
  assign cgp_core_031 = input_a[0] ^ input_b[1];
  assign cgp_core_032 = input_e[2] ^ input_b[1];
  assign cgp_core_033 = input_d[1] & input_d[1];
  assign cgp_core_034 = ~(input_b[0] ^ input_d[1]);
  assign cgp_core_035 = input_d[1] | input_c[1];
  assign cgp_core_036 = input_d[2] ^ input_e[2];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038 = cgp_core_036 ^ cgp_core_035;
  assign cgp_core_039 = cgp_core_036 & cgp_core_035;
  assign cgp_core_040 = cgp_core_037 | cgp_core_039;
  assign cgp_core_043 = input_c[2] | input_d[1];
  assign cgp_core_044 = ~(input_a[2] & input_a[1]);
  assign cgp_core_046 = ~(input_e[0] ^ input_b[2]);
  assign cgp_core_047 = ~(input_e[0] | input_d[2]);
  assign cgp_core_048 = input_c[2] ^ cgp_core_038;
  assign cgp_core_049 = input_c[2] & cgp_core_038;
  assign cgp_core_053 = cgp_core_040 | cgp_core_049;
  assign cgp_core_054 = cgp_core_040 & input_c[2];
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_057 = ~cgp_core_053;
  assign cgp_core_058 = cgp_core_028 & cgp_core_057;
  assign cgp_core_060 = ~(cgp_core_028 ^ cgp_core_053);
  assign cgp_core_061 = cgp_core_060 & cgp_core_056;
  assign cgp_core_062 = ~input_b[2];
  assign cgp_core_064 = cgp_core_026 & cgp_core_061;
  assign cgp_core_065 = ~(input_e[1] | cgp_core_048);
  assign cgp_core_066 = cgp_core_065 & cgp_core_061;
  assign cgp_core_071 = ~(input_d[2] & input_b[1]);
  assign cgp_core_072 = input_c[0] | input_a[1];
  assign cgp_core_074 = ~(input_e[2] & input_a[2]);
  assign cgp_core_076 = input_b[0] ^ input_e[2];
  assign cgp_core_077 = cgp_core_066 | cgp_core_064;
  assign cgp_core_080 = cgp_core_077 | cgp_core_058;

  assign cgp_out[0] = cgp_core_080;
endmodule