module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_069;

  assign cgp_core_014 = input_a[0] ^ input_a[0];
  assign cgp_core_015 = input_d[0] & input_c[0];
  assign cgp_core_016 = input_a[1] ^ input_c[1];
  assign cgp_core_017 = input_a[1] & input_c[1];
  assign cgp_core_018 = ~(input_b[1] | cgp_core_015);
  assign cgp_core_020 = cgp_core_017 | input_d[0];
  assign cgp_core_022 = input_e[0] & input_f[0];
  assign cgp_core_023 = input_e[1] ^ input_a[0];
  assign cgp_core_026 = input_c[1] & cgp_core_022;
  assign cgp_core_027 = input_b[0] | input_a[1];
  assign cgp_core_028_not = ~input_c[1];
  assign cgp_core_032 = input_d[1] ^ input_d[0];
  assign cgp_core_034 = input_e[1] | input_d[0];
  assign cgp_core_035 = input_e[0] ^ cgp_core_034;
  assign cgp_core_037 = input_d[0] | cgp_core_028_not;
  assign cgp_core_038 = input_f[0] & input_c[1];
  assign cgp_core_039 = ~input_f[0];
  assign cgp_core_040 = cgp_core_018 & cgp_core_032;
  assign cgp_core_041 = cgp_core_039 ^ cgp_core_038;
  assign cgp_core_042 = cgp_core_039 & cgp_core_038;
  assign cgp_core_043 = input_a[0] | cgp_core_042;
  assign cgp_core_044 = cgp_core_020 ^ cgp_core_035;
  assign cgp_core_046 = input_f[1] ^ input_e[0];
  assign cgp_core_053 = ~input_e[1];
  assign cgp_core_055 = cgp_core_046 & input_a[0];
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_061 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_062 = cgp_core_061 & input_f[0];
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_064 = ~(input_d[0] & cgp_core_063);
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066 = ~(input_a[0] ^ input_b[0]);
  assign cgp_core_069 = input_d[0] | input_c[0];

  assign cgp_out[0] = 1'b1;
endmodule