module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016_not;
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068_not;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_016_not = ~input_g[1];
  assign cgp_core_017_not = ~input_f[1];
  assign cgp_core_018 = input_e[0] | input_g[1];
  assign cgp_core_023 = ~input_g[0];
  assign cgp_core_026 = input_f[1] & input_a[1];
  assign cgp_core_029 = ~(input_b[1] & input_g[1]);
  assign cgp_core_030 = ~(input_f[1] ^ input_c[0]);
  assign cgp_core_031 = input_d[0] & input_d[1];
  assign cgp_core_032 = ~input_d[0];
  assign cgp_core_034 = ~(input_e[0] & input_c[0]);
  assign cgp_core_035 = ~(input_c[1] & input_b[1]);
  assign cgp_core_036 = ~(input_f[1] ^ input_c[0]);
  assign cgp_core_037 = ~input_a[1];
  assign cgp_core_040 = input_b[1] & input_b[1];
  assign cgp_core_041 = ~input_g[1];
  assign cgp_core_043 = ~(input_f[1] | input_e[1]);
  assign cgp_core_046 = ~(input_d[0] & input_d[1]);
  assign cgp_core_049 = ~(input_a[1] ^ input_d[1]);
  assign cgp_core_053 = ~(input_c[0] ^ input_f[1]);
  assign cgp_core_054 = input_d[0] & input_f[1];
  assign cgp_core_055 = input_e[1] | input_g[0];
  assign cgp_core_056 = input_f[1] ^ input_c[1];
  assign cgp_core_059 = input_f[1] & input_f[1];
  assign cgp_core_061 = ~(input_e[0] ^ input_a[1]);
  assign cgp_core_062 = ~(input_g[1] | input_d[0]);
  assign cgp_core_064 = ~(input_g[1] ^ input_f[0]);
  assign cgp_core_065 = input_f[1] | input_g[0];
  assign cgp_core_066 = ~input_g[0];
  assign cgp_core_068_not = ~input_b[0];
  assign cgp_core_069 = ~(input_d[0] ^ input_d[1]);
  assign cgp_core_070 = ~(input_e[1] & input_b[0]);
  assign cgp_core_073 = ~(input_f[0] & input_e[1]);
  assign cgp_core_075 = ~input_c[1];
  assign cgp_core_076 = input_d[1] | input_c[1];
  assign cgp_core_077 = input_e[1] & input_c[0];
  assign cgp_core_079 = cgp_core_076 | input_g[1];

  assign cgp_out[0] = cgp_core_079;
endmodule