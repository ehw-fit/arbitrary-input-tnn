module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_039_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_062_not;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088_not;
  wire cgp_core_090;

  assign cgp_core_017 = ~(input_a[11] & input_a[8]);
  assign cgp_core_019 = input_a[6] ^ input_a[10];
  assign cgp_core_021 = input_a[6] ^ input_a[7];
  assign cgp_core_022 = ~(input_a[2] | input_a[5]);
  assign cgp_core_024 = input_a[10] & input_a[6];
  assign cgp_core_025 = ~(input_a[7] & input_a[6]);
  assign cgp_core_026 = ~(input_a[3] & input_a[7]);
  assign cgp_core_029 = ~(input_a[0] & input_a[10]);
  assign cgp_core_030 = input_a[9] & input_a[0];
  assign cgp_core_033 = ~(input_a[4] ^ input_a[10]);
  assign cgp_core_034 = input_a[2] ^ input_a[3];
  assign cgp_core_037 = ~input_a[11];
  assign cgp_core_039_not = ~input_a[13];
  assign cgp_core_040 = input_a[4] & input_a[6];
  assign cgp_core_041 = ~(input_a[6] & input_a[7]);
  assign cgp_core_043 = ~(input_a[8] ^ input_a[7]);
  assign cgp_core_045 = ~(input_a[6] ^ input_a[6]);
  assign cgp_core_046 = ~(input_a[5] & input_a[11]);
  assign cgp_core_049 = input_a[1] & input_a[8];
  assign cgp_core_051 = ~(input_a[10] ^ input_a[1]);
  assign cgp_core_053 = input_a[9] | input_a[5];
  assign cgp_core_057 = input_a[8] ^ input_a[4];
  assign cgp_core_058 = input_a[4] ^ input_a[6];
  assign cgp_core_062_not = ~input_a[11];
  assign cgp_core_063 = ~(input_a[3] ^ input_a[0]);
  assign cgp_core_064 = ~cgp_core_049;
  assign cgp_core_065 = input_a[4] & input_a[11];
  assign cgp_core_066 = ~input_a[8];
  assign cgp_core_067 = input_a[6] | input_a[11];
  assign cgp_core_069 = ~input_a[11];
  assign cgp_core_070 = input_a[4] | input_a[1];
  assign cgp_core_071 = ~(input_a[11] ^ input_a[11]);
  assign cgp_core_073 = ~input_a[3];
  assign cgp_core_074_not = ~input_a[8];
  assign cgp_core_075 = input_a[2] | input_a[9];
  assign cgp_core_076 = ~input_a[10];
  assign cgp_core_078 = ~(input_a[3] & input_a[4]);
  assign cgp_core_079 = input_a[13] | input_a[8];
  assign cgp_core_082 = input_a[2] ^ input_a[7];
  assign cgp_core_084 = input_a[13] | input_a[13];
  assign cgp_core_085 = ~input_a[12];
  assign cgp_core_087 = ~(input_a[9] & input_a[6]);
  assign cgp_core_088_not = ~input_a[1];
  assign cgp_core_090 = input_a[0] & input_a[10];

  assign cgp_out[0] = input_a[13];
  assign cgp_out[1] = cgp_core_064;
  assign cgp_out[2] = cgp_core_064;
  assign cgp_out[3] = cgp_core_049;
endmodule