module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047_not;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073_not;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086_not;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092_not;
  wire cgp_core_093;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100_not;
  wire cgp_core_101;
  wire cgp_core_102;
  wire cgp_core_103;
  wire cgp_core_105;

  assign cgp_core_021 = ~(input_g[0] ^ input_c[1]);
  assign cgp_core_024 = ~(input_d[1] | cgp_core_021);
  assign cgp_core_026 = input_f[1] ^ input_d[1];
  assign cgp_core_027 = input_b[1] ^ input_i[1];
  assign cgp_core_028 = input_e[0] & input_c[1];
  assign cgp_core_030 = input_i[0] & input_e[0];
  assign cgp_core_032 = input_f[0] ^ cgp_core_028;
  assign cgp_core_034 = ~(input_b[0] ^ input_a[1]);
  assign cgp_core_036 = ~(input_a[1] | input_h[0]);
  assign cgp_core_037 = ~input_h[1];
  assign cgp_core_038 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_039 = ~(input_h[0] | input_c[0]);
  assign cgp_core_040 = ~(input_e[1] & cgp_core_037);
  assign cgp_core_041 = ~(input_e[0] & input_h[0]);
  assign cgp_core_045 = ~(input_c[0] & input_e[1]);
  assign cgp_core_046 = ~(input_d[0] & input_d[1]);
  assign cgp_core_047_not = ~input_b[0];
  assign cgp_core_050 = input_e[1] | input_b[0];
  assign cgp_core_051 = cgp_core_041 & input_b[0];
  assign cgp_core_052 = input_a[0] & input_e[0];
  assign cgp_core_054 = ~(input_g[1] ^ input_f[0]);
  assign cgp_core_055 = input_f[1] | input_g[0];
  assign cgp_core_056 = input_d[1] ^ input_a[1];
  assign cgp_core_057 = input_c[1] | input_i[0];
  assign cgp_core_060 = ~input_g[1];
  assign cgp_core_061 = ~(input_d[0] | input_c[0]);
  assign cgp_core_062 = input_d[1] ^ input_d[1];
  assign cgp_core_066 = input_c[0] ^ input_e[0];
  assign cgp_core_068 = input_h[0] ^ input_b[0];
  assign cgp_core_069 = input_i[1] & input_h[1];
  assign cgp_core_071 = ~input_g[0];
  assign cgp_core_072 = ~(input_h[1] & input_c[0]);
  assign cgp_core_073_not = ~input_c[0];
  assign cgp_core_076 = input_g[1] & input_c[0];
  assign cgp_core_078 = ~(input_h[0] & input_h[0]);
  assign cgp_core_079 = ~(input_i[1] & input_g[0]);
  assign cgp_core_081 = ~input_b[1];
  assign cgp_core_082 = input_c[0] | input_c[1];
  assign cgp_core_084 = ~(input_h[1] & input_e[1]);
  assign cgp_core_085 = input_e[0] & input_f[0];
  assign cgp_core_086_not = ~input_a[1];
  assign cgp_core_088 = ~(input_d[1] & input_b[1]);
  assign cgp_core_090 = input_g[1] ^ input_e[1];
  assign cgp_core_091 = input_e[0] ^ input_f[0];
  assign cgp_core_092_not = ~input_b[1];
  assign cgp_core_093 = ~(input_d[1] ^ cgp_core_092_not);
  assign cgp_core_096 = ~(input_d[1] ^ input_f[0]);
  assign cgp_core_097 = ~input_e[1];
  assign cgp_core_098 = input_h[1] ^ input_c[1];
  assign cgp_core_099 = input_a[1] | input_c[0];
  assign cgp_core_100_not = ~input_b[1];
  assign cgp_core_101 = input_d[1] & cgp_core_096;
  assign cgp_core_102 = ~(input_b[1] & cgp_core_068);
  assign cgp_core_103 = ~(input_f[1] & input_c[1]);
  assign cgp_core_105 = ~(input_d[0] & cgp_core_068);

  assign cgp_out[0] = 1'b0;
endmodule