module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_050;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_018 = ~(input_c[2] ^ input_c[0]);
  assign cgp_core_019 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_020 = input_a[1] ^ input_c[1];
  assign cgp_core_021 = input_a[2] & cgp_core_018;
  assign cgp_core_022 = ~input_c[1];
  assign cgp_core_025 = input_b[2] ^ input_c[2];
  assign cgp_core_027 = input_c[2] ^ input_d[2];
  assign cgp_core_028 = ~input_c[2];
  assign cgp_core_031 = input_e[0] ^ input_a[2];
  assign cgp_core_032 = input_d[1] ^ input_b[0];
  assign cgp_core_033 = input_e[2] ^ input_d[2];
  assign cgp_core_034 = cgp_core_031 & input_c[0];
  assign cgp_core_037 = input_d[2] & input_d[0];
  assign cgp_core_038 = ~input_b[0];
  assign cgp_core_041_not = ~input_d[0];
  assign cgp_core_042 = ~(input_b[0] | input_c[2]);
  assign cgp_core_043 = input_a[0] ^ input_d[0];
  assign cgp_core_044 = input_a[2] & input_d[2];
  assign cgp_core_045 = input_c[1] ^ input_d[1];
  assign cgp_core_046 = ~(cgp_core_043 & input_a[1]);
  assign cgp_core_050 = ~(input_d[0] | input_d[2]);
  assign cgp_core_056 = input_e[2] ^ input_e[0];
  assign cgp_core_058 = ~(input_d[1] | input_b[1]);
  assign cgp_core_060 = ~input_b[1];
  assign cgp_core_061 = input_a[1] ^ input_b[1];
  assign cgp_core_063 = cgp_core_050 & input_b[1];
  assign cgp_core_066 = ~(input_d[1] ^ cgp_core_050);
  assign cgp_core_068 = ~(cgp_core_045 ^ input_c[2]);
  assign cgp_core_069 = input_a[1] & input_e[1];
  assign cgp_core_071 = ~(input_b[2] | cgp_core_045);
  assign cgp_core_072 = ~(input_a[2] & input_e[1]);
  assign cgp_core_073 = input_c[2] ^ input_d[2];
  assign cgp_core_076 = ~input_e[0];
  assign cgp_core_077 = input_d[2] & cgp_core_072;
  assign cgp_core_078 = ~(input_d[1] | input_c[0]);

  assign cgp_out[0] = 1'b0;
endmodule