module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017 = input_b[2] & input_e[2];
  assign cgp_core_018 = ~(input_d[0] & input_e[0]);
  assign cgp_core_019 = ~input_a[2];
  assign cgp_core_020 = input_e[1] & input_c[1];
  assign cgp_core_024 = input_c[2] | input_e[2];
  assign cgp_core_025 = input_c[2] & input_e[2];
  assign cgp_core_026 = input_e[2] | cgp_core_020;
  assign cgp_core_027 = cgp_core_024 & cgp_core_020;
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_029 = ~(input_e[1] & input_d[0]);
  assign cgp_core_033 = ~(input_e[0] & input_d[2]);
  assign cgp_core_034 = ~input_b[1];
  assign cgp_core_035 = ~(input_d[0] | input_d[2]);
  assign cgp_core_036 = input_b[2] | cgp_core_026;
  assign cgp_core_038 = ~input_d[2];
  assign cgp_core_040 = input_c[2] | cgp_core_036;
  assign cgp_core_041 = input_a[2] | cgp_core_040;
  assign cgp_core_043 = input_c[1] & input_c[1];
  assign cgp_core_044 = ~(input_c[1] | input_b[2]);
  assign cgp_core_045 = input_d[0] | input_d[2];
  assign cgp_core_047 = ~(input_c[0] & input_a[0]);
  assign cgp_core_049 = ~(input_d[2] & input_c[0]);
  assign cgp_core_050 = ~(input_a[0] | input_c[1]);
  assign cgp_core_053 = ~(input_b[0] | input_d[2]);
  assign cgp_core_055 = ~(input_b[0] ^ input_e[2]);
  assign cgp_core_056 = ~input_a[2];
  assign cgp_core_057 = cgp_core_041 & cgp_core_056;
  assign cgp_core_059 = ~input_a[2];
  assign cgp_core_061 = ~(input_d[1] | input_d[1]);
  assign cgp_core_063 = cgp_core_038 & input_b[2];
  assign cgp_core_064 = ~input_b[0];
  assign cgp_core_066 = ~(input_e[0] | input_b[0]);
  assign cgp_core_068 = ~(input_a[0] & input_e[0]);
  assign cgp_core_070 = input_e[1] & input_a[0];
  assign cgp_core_071 = ~(input_d[2] | input_b[0]);
  assign cgp_core_074 = ~(input_c[2] & input_b[2]);
  assign cgp_core_075 = ~input_e[2];
  assign cgp_core_079 = cgp_core_057 | cgp_core_028;
  assign cgp_core_080 = cgp_core_063 | cgp_core_079;

  assign cgp_out[0] = cgp_core_080;
endmodule