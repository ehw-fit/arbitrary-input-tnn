module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031_not;
  wire cgp_core_032;
  wire cgp_core_035_not;
  wire cgp_core_037;
  wire cgp_core_038_not;
  wire cgp_core_039_not;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_053;

  assign cgp_core_012 = input_a[1] | input_e[0];
  assign cgp_core_013 = ~(input_b[0] & input_e[1]);
  assign cgp_core_014 = ~(input_a[1] & input_b[0]);
  assign cgp_core_017 = input_a[1] & input_c[1];
  assign cgp_core_018 = input_e[1] | input_e[1];
  assign cgp_core_019_not = ~input_b[0];
  assign cgp_core_022 = ~(input_b[1] & input_e[0]);
  assign cgp_core_023 = input_e[1] ^ input_a[0];
  assign cgp_core_025 = ~(input_a[1] | input_c[1]);
  assign cgp_core_028 = ~(input_b[0] ^ input_e[1]);
  assign cgp_core_030 = ~(input_c[0] ^ input_d[1]);
  assign cgp_core_031_not = ~input_e[1];
  assign cgp_core_032 = ~(input_a[1] & input_e[1]);
  assign cgp_core_035_not = ~input_c[0];
  assign cgp_core_037 = input_e[0] | input_a[1];
  assign cgp_core_038_not = ~input_e[0];
  assign cgp_core_039_not = ~input_b[0];
  assign cgp_core_040 = ~(input_a[1] | input_c[0]);
  assign cgp_core_042 = ~(input_b[0] | input_e[0]);
  assign cgp_core_045 = ~input_d[1];
  assign cgp_core_046 = ~input_c[0];
  assign cgp_core_047 = input_d[0] ^ input_c[0];
  assign cgp_core_048 = input_c[1] | input_e[0];
  assign cgp_core_053 = input_c[0] | input_d[0];

  assign cgp_out[0] = cgp_core_025;
endmodule