module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065_not;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_072_not;
  wire cgp_core_073;
  wire cgp_core_078;

  assign cgp_core_018 = input_e[0] ^ input_d[2];
  assign cgp_core_019 = input_e[0] | input_b[1];
  assign cgp_core_020 = ~(input_c[2] ^ input_b[2]);
  assign cgp_core_021 = ~(input_d[0] & input_c[1]);
  assign cgp_core_022 = ~input_b[0];
  assign cgp_core_023 = ~(input_a[0] ^ input_c[2]);
  assign cgp_core_024 = ~(input_d[2] & input_a[2]);
  assign cgp_core_025 = input_c[1] | input_e[0];
  assign cgp_core_026 = ~(input_b[1] & input_a[0]);
  assign cgp_core_028 = input_d[1] ^ input_a[0];
  assign cgp_core_029 = input_d[1] ^ input_e[1];
  assign cgp_core_030 = input_a[1] ^ input_c[1];
  assign cgp_core_032 = ~(input_a[0] ^ input_e[2]);
  assign cgp_core_033 = input_b[0] ^ input_a[2];
  assign cgp_core_035 = ~(input_e[2] | input_b[0]);
  assign cgp_core_037 = ~(input_b[0] | input_d[1]);
  assign cgp_core_039 = ~(input_d[1] ^ input_d[1]);
  assign cgp_core_041 = ~(input_b[2] | input_d[0]);
  assign cgp_core_042 = input_e[1] | input_b[0];
  assign cgp_core_043 = ~(input_b[1] & input_d[2]);
  assign cgp_core_044 = ~input_c[0];
  assign cgp_core_048 = ~(input_d[0] | input_c[2]);
  assign cgp_core_049 = input_e[1] ^ input_b[2];
  assign cgp_core_052 = input_c[2] ^ input_d[2];
  assign cgp_core_053 = ~(input_c[1] & input_d[2]);
  assign cgp_core_055 = ~input_e[1];
  assign cgp_core_058 = ~(input_c[2] | input_d[0]);
  assign cgp_core_060 = ~(input_d[1] & input_b[0]);
  assign cgp_core_061 = input_d[0] ^ input_a[0];
  assign cgp_core_063 = input_e[2] ^ input_b[2];
  assign cgp_core_064 = input_b[0] & input_c[1];
  assign cgp_core_065_not = ~input_a[2];
  assign cgp_core_066 = ~input_d[1];
  assign cgp_core_068 = ~input_a[0];
  assign cgp_core_069 = ~input_e[0];
  assign cgp_core_072_not = ~input_a[2];
  assign cgp_core_073 = ~(input_a[2] ^ input_e[0]);
  assign cgp_core_078 = ~(input_a[2] & input_c[0]);

  assign cgp_out[0] = cgp_core_024;
endmodule