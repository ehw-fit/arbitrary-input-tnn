module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_027;
  wire cgp_core_031_not;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046_not;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_078_not;
  wire cgp_core_079;
  wire cgp_core_082;

  assign cgp_core_016 = input_a[0] ^ input_c[0];
  assign cgp_core_017 = input_a[0] & input_c[0];
  assign cgp_core_019 = ~(input_c[1] & input_c[0]);
  assign cgp_core_021 = input_c[0] & input_d[0];
  assign cgp_core_024 = ~input_e[0];
  assign cgp_core_025_not = ~input_g[1];
  assign cgp_core_027 = cgp_core_025_not ^ cgp_core_024;
  assign cgp_core_031_not = ~input_g[1];
  assign cgp_core_032 = ~(input_b[1] & input_f[0]);
  assign cgp_core_033 = input_e[1] & cgp_core_027;
  assign cgp_core_034 = input_a[0] ^ input_b[1];
  assign cgp_core_037_not = ~input_d[1];
  assign cgp_core_040 = input_g[1] & input_a[0];
  assign cgp_core_041 = input_b[1] ^ cgp_core_034;
  assign cgp_core_042 = ~(input_c[0] ^ cgp_core_034);
  assign cgp_core_043 = input_c[0] ^ input_b[1];
  assign cgp_core_046_not = ~cgp_core_037_not;
  assign cgp_core_048 = input_d[0] ^ input_c[0];
  assign cgp_core_050 = input_e[1] & input_b[0];
  assign cgp_core_053 = input_b[1] ^ input_f[0];
  assign cgp_core_055 = input_b[1] ^ input_d[1];
  assign cgp_core_060 = ~input_c[1];
  assign cgp_core_064 = input_b[1] & input_c[1];
  assign cgp_core_066 = cgp_core_048 & input_a[1];
  assign cgp_core_067 = ~(input_c[0] | input_g[0]);
  assign cgp_core_071 = ~(input_d[1] | input_a[1]);
  assign cgp_core_072 = cgp_core_043 | input_f[1];
  assign cgp_core_073 = input_b[1] ^ input_b[0];
  assign cgp_core_074 = input_a[1] & input_b[0];
  assign cgp_core_078_not = ~cgp_core_073;
  assign cgp_core_079 = ~(input_e[0] | input_g[1]);
  assign cgp_core_082 = ~(input_g[1] | input_f[1]);

  assign cgp_out[0] = 1'b1;
endmodule