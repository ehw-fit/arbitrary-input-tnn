module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012_not;
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_012_not = ~input_c[0];
  assign cgp_core_014 = ~(input_e[0] & input_b[1]);
  assign cgp_core_016 = input_e[0] | input_a[0];
  assign cgp_core_020 = ~input_d[0];
  assign cgp_core_023 = ~(input_d[1] ^ input_c[1]);
  assign cgp_core_024 = ~input_e[0];
  assign cgp_core_025 = input_e[1] | input_c[1];
  assign cgp_core_029 = input_e[1] ^ input_a[0];
  assign cgp_core_031 = ~(input_b[0] & input_b[1]);
  assign cgp_core_032 = input_a[0] ^ input_b[0];
  assign cgp_core_033 = cgp_core_025 | input_a[1];
  assign cgp_core_034 = cgp_core_025 & input_a[1];
  assign cgp_core_035 = ~input_a[0];
  assign cgp_core_036 = ~cgp_core_034;
  assign cgp_core_037 = ~cgp_core_033;
  assign cgp_core_041 = input_d[1] & cgp_core_036;
  assign cgp_core_043 = ~input_d[0];
  assign cgp_core_045 = input_d[0] ^ input_d[1];
  assign cgp_core_051 = input_b[1] & cgp_core_041;
  assign cgp_core_052 = ~input_e[0];
  assign cgp_core_053 = cgp_core_037 | cgp_core_051;
  assign cgp_core_054 = ~input_d[0];

  assign cgp_out[0] = cgp_core_053;
endmodule