module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016_not;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_015 = ~input_b[1];
  assign cgp_core_016_not = ~input_c[0];
  assign cgp_core_020 = input_e[1] | input_e[0];
  assign cgp_core_021 = ~(input_e[0] | input_f[1]);
  assign cgp_core_023 = ~input_a[1];
  assign cgp_core_025 = input_f[0] ^ input_e[0];
  assign cgp_core_026 = ~(input_e[1] | input_e[0]);
  assign cgp_core_027 = input_a[0] & input_a[0];
  assign cgp_core_028 = input_c[1] ^ input_c[0];
  assign cgp_core_030 = ~(input_c[0] & input_a[1]);
  assign cgp_core_033 = ~input_d[0];
  assign cgp_core_034 = input_f[0] ^ input_f[0];
  assign cgp_core_035 = ~(input_f[1] | input_d[1]);
  assign cgp_core_036 = input_b[1] ^ input_b[0];
  assign cgp_core_037 = input_e[1] | input_c[0];
  assign cgp_core_040 = input_f[0] & input_c[1];
  assign cgp_core_043 = input_d[1] ^ input_f[0];
  assign cgp_core_044 = cgp_core_020 | input_a[0];
  assign cgp_core_045 = ~(input_c[0] & input_f[1]);
  assign cgp_core_047 = input_b[0] ^ input_d[1];
  assign cgp_core_049_not = ~input_c[1];
  assign cgp_core_050 = ~input_c[1];
  assign cgp_core_051 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_056 = ~(input_d[0] | input_b[1]);
  assign cgp_core_058 = input_b[0] ^ input_c[1];
  assign cgp_core_059 = ~(input_c[1] & input_d[0]);
  assign cgp_core_060 = input_c[1] & input_f[0];
  assign cgp_core_061 = input_e[1] | input_f[1];
  assign cgp_core_062 = ~input_b[1];
  assign cgp_core_063 = input_d[0] ^ input_f[1];
  assign cgp_core_066 = input_f[1] ^ input_e[1];
  assign cgp_core_067 = ~(input_a[0] & input_f[1]);
  assign cgp_core_068 = input_a[1] | cgp_core_044;
  assign cgp_core_069 = input_f[1] | cgp_core_068;
  assign cgp_core_070 = input_d[1] | input_d[0];
  assign cgp_core_071 = input_c[1] | cgp_core_070;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;

  assign cgp_out[0] = cgp_core_072;
endmodule