module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019_not;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_066;

  assign cgp_core_017 = ~input_a[1];
  assign cgp_core_019_not = ~input_b[0];
  assign cgp_core_020 = ~(cgp_core_017 & input_e[0]);
  assign cgp_core_021 = input_b[0] & input_e[1];
  assign cgp_core_022 = ~(input_b[0] | input_c[0]);
  assign cgp_core_023 = input_b[1] & input_d[1];
  assign cgp_core_024_not = ~input_a[0];
  assign cgp_core_025 = input_c[0] ^ cgp_core_022;
  assign cgp_core_026 = input_b[0] | input_c[0];
  assign cgp_core_027 = ~(input_e[0] & cgp_core_026);
  assign cgp_core_030 = input_a[1] ^ input_a[1];
  assign cgp_core_031 = ~input_e[1];
  assign cgp_core_033 = input_e[1] & input_b[0];
  assign cgp_core_035 = input_c[0] | input_b[0];
  assign cgp_core_037 = ~(input_c[0] & input_f[1]);
  assign cgp_core_039 = ~(input_c[0] ^ input_c[0]);
  assign cgp_core_040 = ~cgp_core_037;
  assign cgp_core_041 = ~(input_a[1] & cgp_core_040);
  assign cgp_core_043 = cgp_core_027 & input_f[1];
  assign cgp_core_044 = input_c[0] ^ cgp_core_041;
  assign cgp_core_047 = input_a[1] ^ input_a[0];
  assign cgp_core_048 = ~input_a[0];
  assign cgp_core_055 = input_b[1] | input_e[0];
  assign cgp_core_057 = ~(input_e[1] | cgp_core_039);
  assign cgp_core_066 = input_a[0] | input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule