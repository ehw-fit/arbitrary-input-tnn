module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061_not;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068_not;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_021 = ~(input_b[0] ^ input_a[0]);
  assign cgp_core_022 = ~(input_b[2] | input_e[1]);
  assign cgp_core_023 = ~(input_b[0] ^ input_b[1]);
  assign cgp_core_024 = ~(input_e[1] ^ input_c[1]);
  assign cgp_core_025 = input_f[0] & input_a[0];
  assign cgp_core_026_not = ~input_c[0];
  assign cgp_core_028 = input_c[2] & input_e[2];
  assign cgp_core_029 = ~(input_d[2] ^ input_a[1]);
  assign cgp_core_030 = input_b[2] | input_d[0];
  assign cgp_core_034 = ~(input_d[0] & input_e[0]);
  assign cgp_core_035 = ~(input_e[0] ^ input_e[2]);
  assign cgp_core_038 = input_a[0] & input_d[1];
  assign cgp_core_039 = input_b[2] & input_d[0];
  assign cgp_core_041 = ~input_d[2];
  assign cgp_core_042 = input_e[0] | input_b[0];
  assign cgp_core_044 = cgp_core_028 | input_a[2];
  assign cgp_core_045 = cgp_core_028 & input_a[2];
  assign cgp_core_046 = ~(input_b[1] ^ input_e[1]);
  assign cgp_core_047 = ~(input_e[0] | input_f[2]);
  assign cgp_core_049 = input_d[2] | input_c[2];
  assign cgp_core_051 = input_b[0] | input_d[0];
  assign cgp_core_053 = ~(input_f[1] | input_f[0]);
  assign cgp_core_055 = input_b[2] | input_b[0];
  assign cgp_core_056 = ~input_e[0];
  assign cgp_core_057 = ~(input_d[1] ^ input_d[0]);
  assign cgp_core_058 = ~input_a[2];
  assign cgp_core_059 = input_c[1] & input_b[1];
  assign cgp_core_060 = input_c[2] & input_e[1];
  assign cgp_core_061_not = ~input_e[1];
  assign cgp_core_064 = ~(input_b[1] & input_a[1]);
  assign cgp_core_065 = ~(input_e[2] | input_c[1]);
  assign cgp_core_066 = input_b[2] ^ input_c[2];
  assign cgp_core_068_not = ~input_f[2];
  assign cgp_core_069 = input_b[2] | input_d[2];
  assign cgp_core_070 = input_d[2] | input_b[2];
  assign cgp_core_071 = input_f[2] & cgp_core_069;
  assign cgp_core_074_not = ~cgp_core_071;
  assign cgp_core_075 = input_e[1] & input_a[2];
  assign cgp_core_077 = cgp_core_044 & cgp_core_074_not;
  assign cgp_core_078 = ~(input_f[2] | cgp_core_070);
  assign cgp_core_080 = ~input_e[1];
  assign cgp_core_086 = ~(input_b[2] & input_b[1]);
  assign cgp_core_087 = ~(input_b[1] & input_c[1]);
  assign cgp_core_089 = ~(input_f[2] ^ input_a[2]);
  assign cgp_core_090 = ~(input_a[1] | input_f[2]);
  assign cgp_core_091 = ~(input_d[0] & input_f[2]);
  assign cgp_core_093 = ~(input_f[0] | input_f[2]);
  assign cgp_core_098 = cgp_core_077 | cgp_core_045;
  assign cgp_core_099 = cgp_core_078 | cgp_core_098;

  assign cgp_out[0] = cgp_core_099;
endmodule