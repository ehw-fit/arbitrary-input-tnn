module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_030;
  wire cgp_core_031_not;
  wire cgp_core_036;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046_not;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_018 = input_b[2] & input_b[0];
  assign cgp_core_019 = input_c[1] & input_d[0];
  assign cgp_core_020 = ~(input_c[1] ^ input_e[1]);
  assign cgp_core_022 = ~(input_d[1] & input_e[1]);
  assign cgp_core_025 = input_b[0] & input_e[2];
  assign cgp_core_030 = input_b[0] & input_e[0];
  assign cgp_core_031_not = ~input_a[1];
  assign cgp_core_036 = ~(input_e[1] | input_d[2]);
  assign cgp_core_041_not = ~input_e[1];
  assign cgp_core_042 = ~(input_b[2] & input_e[1]);
  assign cgp_core_043 = input_d[0] ^ input_b[0];
  assign cgp_core_044 = input_a[0] | input_c[1];
  assign cgp_core_045 = input_a[1] & input_d[1];
  assign cgp_core_046_not = ~input_a[1];
  assign cgp_core_047 = cgp_core_045 ^ cgp_core_044;
  assign cgp_core_048 = input_b[2] ^ input_d[1];
  assign cgp_core_050 = input_a[2] ^ input_c[2];
  assign cgp_core_055 = input_c[2] & input_b[2];
  assign cgp_core_056 = ~input_b[0];
  assign cgp_core_057 = input_c[0] & cgp_core_056;
  assign cgp_core_058 = cgp_core_057 & cgp_core_055;
  assign cgp_core_061 = ~(input_e[0] ^ input_c[2]);
  assign cgp_core_062 = input_a[0] & input_c[1];
  assign cgp_core_063 = input_c[1] & input_d[0];
  assign cgp_core_065 = ~input_d[0];
  assign cgp_core_066 = ~(cgp_core_047 ^ cgp_core_047);
  assign cgp_core_067 = input_c[2] & cgp_core_066;
  assign cgp_core_068 = cgp_core_067 & cgp_core_065;
  assign cgp_core_069 = ~(input_d[1] | input_b[1]);
  assign cgp_core_071 = ~cgp_core_043;
  assign cgp_core_076 = input_e[0] | input_a[0];
  assign cgp_core_077 = input_d[2] | cgp_core_076;
  assign cgp_core_078 = input_a[0] | input_c[2];
  assign cgp_core_079 = ~(input_a[1] | input_e[0]);
  assign cgp_core_080 = input_c[1] | input_e[1];

  assign cgp_out[0] = 1'b1;
endmodule