module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_078_not;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_083;

  assign cgp_core_016 = ~(input_a[0] ^ input_a[0]);
  assign cgp_core_018 = ~(input_g[1] & input_b[0]);
  assign cgp_core_019 = input_a[0] & input_b[1];
  assign cgp_core_020 = input_e[0] & input_f[1];
  assign cgp_core_022 = ~(input_g[1] ^ input_e[0]);
  assign cgp_core_024 = ~input_b[0];
  assign cgp_core_025 = input_g[0] | input_g[0];
  assign cgp_core_027 = input_g[0] ^ input_f[0];
  assign cgp_core_029 = input_d[0] | input_c[0];
  assign cgp_core_030 = input_f[1] | input_g[1];
  assign cgp_core_032 = ~input_c[0];
  assign cgp_core_034 = ~(input_b[0] ^ input_e[0]);
  assign cgp_core_036 = input_e[1] & input_d[0];
  assign cgp_core_038 = input_d[0] & input_g[1];
  assign cgp_core_041 = ~input_g[0];
  assign cgp_core_046 = input_e[0] | input_c[0];
  assign cgp_core_048 = input_g[1] | input_e[1];
  assign cgp_core_049_not = ~input_b[1];
  assign cgp_core_050 = ~(input_e[1] | input_b[0]);
  assign cgp_core_051 = ~(input_b[1] & input_g[0]);
  assign cgp_core_052 = input_c[0] | input_b[1];
  assign cgp_core_056 = ~(input_g[1] & input_d[0]);
  assign cgp_core_058 = ~(input_g[0] & input_e[1]);
  assign cgp_core_059 = ~(input_c[1] | input_d[1]);
  assign cgp_core_060 = ~input_f[1];
  assign cgp_core_063 = input_b[1] | input_c[0];
  assign cgp_core_064 = ~(input_c[1] ^ input_g[1]);
  assign cgp_core_067 = ~(input_f[0] | input_e[1]);
  assign cgp_core_068 = input_d[0] | input_a[0];
  assign cgp_core_070 = input_a[0] | input_c[0];
  assign cgp_core_073 = input_g[1] | input_b[0];
  assign cgp_core_076 = input_e[0] ^ input_b[1];
  assign cgp_core_078_not = ~input_b[0];
  assign cgp_core_079 = input_d[1] | cgp_core_048;
  assign cgp_core_080 = input_c[1] | cgp_core_079;
  assign cgp_core_083 = cgp_core_080 | input_a[1];

  assign cgp_out[0] = cgp_core_083;
endmodule