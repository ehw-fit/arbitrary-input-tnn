module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_031_not;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_039;

  assign cgp_core_012 = input_c[1] ^ input_d[1];
  assign cgp_core_013 = input_c[1] & input_d[1];
  assign cgp_core_014 = cgp_core_012 ^ input_c[0];
  assign cgp_core_015 = input_a[1] & input_c[0];
  assign cgp_core_016 = cgp_core_013 | input_a[0];
  assign cgp_core_018 = input_b[0] & input_c[0];
  assign cgp_core_019 = ~(input_b[0] | input_c[0]);
  assign cgp_core_020 = input_a[0] & cgp_core_014;
  assign cgp_core_021 = cgp_core_019 ^ cgp_core_018;
  assign cgp_core_022 = cgp_core_019 & cgp_core_018;
  assign cgp_core_023 = input_c[0] | cgp_core_022;
  assign cgp_core_025 = cgp_core_016 & cgp_core_023;
  assign cgp_core_026 = ~cgp_core_025;
  assign cgp_core_027_not = ~cgp_core_026;
  assign cgp_core_031_not = ~input_d[1];
  assign cgp_core_033 = ~(cgp_core_021 ^ input_a[1]);
  assign cgp_core_035 = ~input_a[0];
  assign cgp_core_039 = input_a[0] & cgp_core_033;

  assign cgp_out[0] = 1'b1;
endmodule