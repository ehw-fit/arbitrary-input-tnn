module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015_not;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_013 = ~(input_d[1] & input_e[0]);
  assign cgp_core_014 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_015_not = ~input_e[1];
  assign cgp_core_017 = ~input_c[1];
  assign cgp_core_019 = input_d[1] & input_d[0];
  assign cgp_core_021 = ~input_a[1];
  assign cgp_core_022 = input_d[0] & input_a[1];
  assign cgp_core_025 = ~(input_d[1] & input_c[1]);
  assign cgp_core_026 = input_b[0] & input_a[0];
  assign cgp_core_027 = ~(input_e[1] ^ input_c[1]);
  assign cgp_core_029 = input_a[0] & input_b[0];
  assign cgp_core_030 = ~input_c[0];
  assign cgp_core_032 = input_e[0] | input_a[0];
  assign cgp_core_033 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_038 = input_e[1] | input_b[1];
  assign cgp_core_040 = ~input_b[0];
  assign cgp_core_042 = ~input_c[0];
  assign cgp_core_043 = input_e[0] & input_c[1];
  assign cgp_core_045 = ~input_a[1];
  assign cgp_core_049 = input_a[1] | input_a[0];
  assign cgp_core_052 = input_c[0] ^ input_d[1];
  assign cgp_core_053 = ~(input_c[0] & input_a[1]);
  assign cgp_core_054 = input_e[0] | input_b[1];

  assign cgp_out[0] = cgp_core_025;
endmodule