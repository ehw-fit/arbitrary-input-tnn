module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016_not;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047_not;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070_not;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;

  assign cgp_core_016_not = ~input_a[13];
  assign cgp_core_018 = ~(input_a[10] & input_a[5]);
  assign cgp_core_019 = ~(input_a[13] & input_a[7]);
  assign cgp_core_020 = ~(input_a[7] & input_a[13]);
  assign cgp_core_022 = ~(input_a[11] ^ input_a[10]);
  assign cgp_core_025_not = ~input_a[10];
  assign cgp_core_026 = input_a[9] & input_a[2];
  assign cgp_core_027 = input_a[3] & input_a[8];
  assign cgp_core_029 = input_a[9] ^ input_a[3];
  assign cgp_core_030 = ~(input_a[7] | input_a[6]);
  assign cgp_core_031 = input_a[10] & input_a[2];
  assign cgp_core_032 = input_a[11] ^ input_a[11];
  assign cgp_core_035_not = ~input_a[2];
  assign cgp_core_037 = ~(input_a[8] & input_a[0]);
  assign cgp_core_038 = input_a[8] & input_a[0];
  assign cgp_core_043 = ~input_a[9];
  assign cgp_core_044 = input_a[7] | input_a[9];
  assign cgp_core_047_not = ~input_a[3];
  assign cgp_core_048 = input_a[7] & input_a[1];
  assign cgp_core_049 = ~(input_a[0] & input_a[12]);
  assign cgp_core_051 = ~(input_a[3] ^ input_a[3]);
  assign cgp_core_054 = ~(input_a[7] & input_a[2]);
  assign cgp_core_055 = input_a[7] ^ input_a[8];
  assign cgp_core_057 = ~input_a[0];
  assign cgp_core_058 = input_a[0] ^ input_a[12];
  assign cgp_core_059 = ~(input_a[8] & input_a[7]);
  assign cgp_core_061 = ~(input_a[5] | input_a[3]);
  assign cgp_core_064 = ~input_a[5];
  assign cgp_core_066 = cgp_core_064 ^ input_a[6];
  assign cgp_core_068 = input_a[0] ^ input_a[10];
  assign cgp_core_070_not = ~input_a[1];
  assign cgp_core_071 = input_a[5] | input_a[6];
  assign cgp_core_072 = ~(input_a[2] | input_a[0]);
  assign cgp_core_073 = ~(input_a[6] ^ input_a[1]);
  assign cgp_core_076 = input_a[6] | input_a[5];
  assign cgp_core_077 = cgp_core_037 & cgp_core_066;
  assign cgp_core_078 = ~(input_a[7] ^ input_a[2]);
  assign cgp_core_079 = input_a[2] ^ input_a[1];
  assign cgp_core_081 = cgp_core_038 ^ cgp_core_071;
  assign cgp_core_082 = cgp_core_038 & cgp_core_071;
  assign cgp_core_083 = cgp_core_081 ^ cgp_core_077;
  assign cgp_core_084 = input_a[5] & input_a[6];
  assign cgp_core_085 = cgp_core_082 | cgp_core_084;
  assign cgp_core_087 = input_a[12] ^ input_a[13];
  assign cgp_core_088 = input_a[9] | input_a[6];
  assign cgp_core_089 = ~input_a[13];

  assign cgp_out[0] = 1'b0;
  assign cgp_out[1] = cgp_core_083;
  assign cgp_out[2] = cgp_core_083;
  assign cgp_out[3] = cgp_core_085;
endmodule