module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061_not;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_071;

  assign cgp_core_014 = input_e[0] ^ input_c[0];
  assign cgp_core_016 = input_a[1] & input_c[1];
  assign cgp_core_017 = input_a[1] & input_c[1];
  assign cgp_core_021 = input_e[0] ^ input_f[0];
  assign cgp_core_022 = input_e[0] & input_f[0];
  assign cgp_core_023 = input_b[1] ^ input_f[1];
  assign cgp_core_024 = input_e[1] & input_f[1];
  assign cgp_core_025 = cgp_core_023 ^ cgp_core_022;
  assign cgp_core_026 = ~(input_f[0] & input_d[1]);
  assign cgp_core_027 = cgp_core_024 | input_d[0];
  assign cgp_core_028 = input_d[0] ^ cgp_core_021;
  assign cgp_core_029 = input_c[0] & input_c[0];
  assign cgp_core_030 = input_d[1] ^ cgp_core_025;
  assign cgp_core_031 = ~(input_e[1] | input_e[1]);
  assign cgp_core_035 = input_f[1] ^ cgp_core_031;
  assign cgp_core_037 = ~(input_c[1] & cgp_core_028);
  assign cgp_core_038 = cgp_core_014 ^ input_b[1];
  assign cgp_core_039_not = ~input_e[1];
  assign cgp_core_041 = cgp_core_039_not ^ cgp_core_038;
  assign cgp_core_042 = input_a[1] & cgp_core_038;
  assign cgp_core_044 = cgp_core_016 ^ cgp_core_035;
  assign cgp_core_045 = ~cgp_core_016;
  assign cgp_core_046 = cgp_core_044 & input_d[1];
  assign cgp_core_047 = ~(cgp_core_044 | input_f[1]);
  assign cgp_core_048 = ~(input_c[1] & input_d[1]);
  assign cgp_core_049_not = ~cgp_core_048;
  assign cgp_core_051 = ~input_d[0];
  assign cgp_core_052 = cgp_core_049_not & input_f[0];
  assign cgp_core_053 = ~cgp_core_049_not;
  assign cgp_core_054 = cgp_core_053 & cgp_core_051;
  assign cgp_core_055 = cgp_core_046 ^ cgp_core_054;
  assign cgp_core_056 = ~cgp_core_046;
  assign cgp_core_057 = input_c[0] & input_e[0];
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_059 = input_c[1] & input_c[1];
  assign cgp_core_060 = input_d[1] & cgp_core_057;
  assign cgp_core_061_not = ~input_f[1];
  assign cgp_core_062 = input_e[0] & input_c[1];
  assign cgp_core_063 = ~input_a[1];
  assign cgp_core_064_not = ~input_c[1];
  assign cgp_core_066 = ~(cgp_core_037 ^ input_b[0]);
  assign cgp_core_067 = input_c[0] & input_d[0];
  assign cgp_core_071 = ~(cgp_core_052 & input_c[1]);

  assign cgp_out[0] = 1'b1;
endmodule