module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_010;
  wire cgp_core_014_not;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027_not;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;

  assign cgp_core_010 = input_c[0] ^ input_d[0];
  assign cgp_core_014_not = ~input_b[1];
  assign cgp_core_017 = input_d[0] & input_c[1];
  assign cgp_core_018 = input_a[1] & input_d[1];
  assign cgp_core_019 = ~(input_b[0] & input_b[1]);
  assign cgp_core_021 = input_b[1] & input_b[1];
  assign cgp_core_024 = ~(input_c[1] | input_a[0]);
  assign cgp_core_025 = input_a[0] & input_b[1];
  assign cgp_core_027_not = ~input_a[1];
  assign cgp_core_028 = ~(input_d[1] & input_d[0]);
  assign cgp_core_030 = ~(input_d[0] & input_c[0]);
  assign cgp_core_031 = input_d[1] | input_a[0];
  assign cgp_core_034 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_036 = ~(input_a[1] & input_b[1]);
  assign cgp_core_037 = input_c[0] ^ input_a[0];
  assign cgp_core_040 = input_c[1] | input_d[1];
  assign cgp_core_042 = input_b[1] | input_c[0];
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;

  assign cgp_out[0] = cgp_core_043;
endmodule