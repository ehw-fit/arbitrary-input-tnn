module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_023;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066_not;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_088;
  wire cgp_core_092;

  assign cgp_core_019 = ~(input_a[1] | input_g[0]);
  assign cgp_core_023 = ~input_b[0];
  assign cgp_core_026_not = ~input_c[1];
  assign cgp_core_027 = ~(input_a[1] & input_h[1]);
  assign cgp_core_032 = ~(input_f[0] | input_h[0]);
  assign cgp_core_035 = ~(input_a[1] | input_h[1]);
  assign cgp_core_036 = input_b[1] & input_e[0];
  assign cgp_core_038 = ~input_f[0];
  assign cgp_core_039 = input_h[1] & input_c[0];
  assign cgp_core_040 = input_f[1] | input_b[0];
  assign cgp_core_041 = ~(input_a[0] | input_h[1]);
  assign cgp_core_044 = ~input_e[1];
  assign cgp_core_045 = input_e[1] ^ input_b[0];
  assign cgp_core_049 = input_g[1] & input_e[1];
  assign cgp_core_050 = ~input_c[0];
  assign cgp_core_051 = input_h[0] & cgp_core_045;
  assign cgp_core_053 = ~(input_b[0] ^ input_f[1]);
  assign cgp_core_054 = input_b[1] | input_c[0];
  assign cgp_core_057 = input_e[1] | input_f[1];
  assign cgp_core_058 = ~input_c[0];
  assign cgp_core_062 = input_c[0] ^ input_h[0];
  assign cgp_core_063 = ~(input_h[0] ^ input_b[1]);
  assign cgp_core_064 = ~input_f[0];
  assign cgp_core_066_not = ~cgp_core_063;
  assign cgp_core_067 = ~(input_e[0] | input_h[0]);
  assign cgp_core_069 = input_e[1] | input_h[1];
  assign cgp_core_073 = ~input_h[0];
  assign cgp_core_075 = input_a[1] & input_d[1];
  assign cgp_core_077 = input_e[1] & input_e[0];
  assign cgp_core_078 = ~(input_f[0] | input_d[1]);
  assign cgp_core_080 = ~input_b[1];
  assign cgp_core_081 = input_g[0] & cgp_core_066_not;
  assign cgp_core_082 = ~(cgp_core_081 & input_g[0]);
  assign cgp_core_084 = cgp_core_027 & input_g[0];
  assign cgp_core_085 = ~(input_e[0] | input_a[0]);
  assign cgp_core_088 = ~(cgp_core_057 | input_d[1]);
  assign cgp_core_092 = input_e[1] & cgp_core_082;

  assign cgp_out[0] = 1'b0;
endmodule