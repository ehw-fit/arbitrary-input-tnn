module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055_not;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075_not;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;

  assign cgp_core_016 = input_a[2] ^ input_a[12];
  assign cgp_core_017 = input_a[0] & input_a[11];
  assign cgp_core_018 = ~input_a[8];
  assign cgp_core_021 = input_a[10] & input_a[10];
  assign cgp_core_023 = ~(input_a[1] | input_a[10]);
  assign cgp_core_025 = ~input_a[3];
  assign cgp_core_029 = ~(input_a[2] & input_a[13]);
  assign cgp_core_030 = ~(input_a[4] | input_a[13]);
  assign cgp_core_033 = input_a[5] & input_a[12];
  assign cgp_core_035 = ~(input_a[4] ^ input_a[1]);
  assign cgp_core_037 = ~input_a[11];
  assign cgp_core_038 = input_a[8] ^ input_a[5];
  assign cgp_core_039 = input_a[2] | input_a[12];
  assign cgp_core_040 = input_a[7] | input_a[7];
  assign cgp_core_041 = ~(input_a[4] ^ input_a[1]);
  assign cgp_core_042_not = ~input_a[6];
  assign cgp_core_043 = input_a[2] | input_a[4];
  assign cgp_core_044 = input_a[4] | input_a[8];
  assign cgp_core_045 = ~(input_a[7] ^ input_a[1]);
  assign cgp_core_046 = ~(input_a[0] & input_a[5]);
  assign cgp_core_048 = ~(input_a[1] | input_a[8]);
  assign cgp_core_052 = ~input_a[0];
  assign cgp_core_054 = input_a[2] | input_a[7];
  assign cgp_core_055_not = ~input_a[6];
  assign cgp_core_057 = ~(input_a[5] | input_a[12]);
  assign cgp_core_059 = ~(input_a[10] | input_a[7]);
  assign cgp_core_060 = ~(input_a[4] & input_a[8]);
  assign cgp_core_065 = ~input_a[1];
  assign cgp_core_067 = input_a[8] & input_a[8];
  assign cgp_core_069 = ~(input_a[4] | input_a[2]);
  assign cgp_core_071 = ~(input_a[0] & input_a[2]);
  assign cgp_core_072 = ~input_a[12];
  assign cgp_core_073 = input_a[8] & input_a[1];
  assign cgp_core_074 = ~(input_a[2] & input_a[9]);
  assign cgp_core_075_not = ~input_a[12];
  assign cgp_core_081 = input_a[2] & input_a[3];
  assign cgp_core_083 = ~cgp_core_081;
  assign cgp_core_084 = ~input_a[1];
  assign cgp_core_085 = ~(input_a[1] ^ input_a[4]);
  assign cgp_core_086 = input_a[13] ^ input_a[7];

  assign cgp_out[0] = input_a[9];
  assign cgp_out[1] = cgp_core_083;
  assign cgp_out[2] = cgp_core_083;
  assign cgp_out[3] = cgp_core_081;
endmodule