module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_071;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_091;
  wire cgp_core_092;

  assign cgp_core_018 = input_e[1] | input_f[1];
  assign cgp_core_020 = input_c[0] ^ input_h[1];
  assign cgp_core_021 = input_d[1] & input_a[0];
  assign cgp_core_022 = input_a[1] ^ input_a[0];
  assign cgp_core_024 = input_h[0] | input_e[1];
  assign cgp_core_026 = ~(input_a[0] ^ input_g[0]);
  assign cgp_core_027 = input_e[0] & input_b[1];
  assign cgp_core_028 = input_f[0] ^ input_f[0];
  assign cgp_core_029_not = ~input_b[1];
  assign cgp_core_032_not = ~input_h[0];
  assign cgp_core_033 = input_c[1] & input_e[1];
  assign cgp_core_034 = input_c[0] ^ input_a[0];
  assign cgp_core_039 = input_f[1] & input_g[0];
  assign cgp_core_040 = input_a[1] & input_e[0];
  assign cgp_core_042 = input_f[1] | input_h[1];
  assign cgp_core_044 = ~(input_f[1] | input_e[1]);
  assign cgp_core_045 = ~(input_e[1] | input_f[0]);
  assign cgp_core_046 = ~(input_c[0] ^ input_g[0]);
  assign cgp_core_047 = cgp_core_044 | input_h[0];
  assign cgp_core_049 = ~(input_h[1] | input_c[1]);
  assign cgp_core_050 = input_d[0] ^ input_g[0];
  assign cgp_core_051 = ~(input_c[1] & cgp_core_045);
  assign cgp_core_052 = ~(cgp_core_050 & input_e[0]);
  assign cgp_core_055 = ~cgp_core_047;
  assign cgp_core_059 = ~(input_d[1] & input_c[0]);
  assign cgp_core_060 = ~input_f[1];
  assign cgp_core_064 = ~input_f[0];
  assign cgp_core_066 = cgp_core_064 | input_d[1];
  assign cgp_core_067 = input_h[1] | input_d[1];
  assign cgp_core_071 = ~input_d[0];
  assign cgp_core_080 = ~input_a[1];
  assign cgp_core_081 = ~(input_e[0] ^ cgp_core_066);
  assign cgp_core_082 = ~(input_a[1] ^ input_d[1]);
  assign cgp_core_083 = ~(input_d[0] & input_b[1]);
  assign cgp_core_084 = input_e[0] & input_d[1];
  assign cgp_core_085 = input_h[0] & input_d[0];
  assign cgp_core_087 = input_d[1] | cgp_core_082;
  assign cgp_core_091 = ~input_b[1];
  assign cgp_core_092 = input_d[1] & input_e[0];

  assign cgp_out[0] = 1'b0;
endmodule