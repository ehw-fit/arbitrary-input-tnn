module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_038;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_068;
  wire cgp_core_071;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_091;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_099;
  wire cgp_core_101;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_107;

  assign cgp_core_020 = input_i[0] & input_h[0];
  assign cgp_core_022 = ~input_a[1];
  assign cgp_core_023 = ~(input_a[0] ^ input_i[1]);
  assign cgp_core_024 = ~(cgp_core_022 ^ input_i[0]);
  assign cgp_core_026 = input_a[0] | input_a[1];
  assign cgp_core_027 = input_f[0] | input_d[0];
  assign cgp_core_028 = input_h[1] ^ input_b[0];
  assign cgp_core_030 = ~input_c[1];
  assign cgp_core_031 = input_i[0] | input_c[1];
  assign cgp_core_032_not = ~input_h[0];
  assign cgp_core_033 = input_a[0] ^ input_b[0];
  assign cgp_core_038 = input_h[0] & input_f[1];
  assign cgp_core_041_not = ~input_g[0];
  assign cgp_core_042 = input_e[1] ^ input_e[1];
  assign cgp_core_049 = input_f[1] & input_e[0];
  assign cgp_core_050 = cgp_core_042 ^ input_a[1];
  assign cgp_core_052 = ~(input_i[1] & input_g[1]);
  assign cgp_core_053 = ~input_g[1];
  assign cgp_core_054 = ~(input_h[1] | input_f[0]);
  assign cgp_core_055 = input_a[0] & input_g[1];
  assign cgp_core_056 = ~(cgp_core_054 ^ input_c[0]);
  assign cgp_core_058 = ~(input_b[1] ^ input_b[0]);
  assign cgp_core_059 = input_a[0] & input_a[0];
  assign cgp_core_061 = input_c[1] & input_h[0];
  assign cgp_core_068 = input_b[0] ^ input_f[0];
  assign cgp_core_071 = input_e[1] | input_d[0];
  assign cgp_core_075 = ~input_a[0];
  assign cgp_core_078 = ~(input_i[0] & input_b[1]);
  assign cgp_core_079 = ~input_d[1];
  assign cgp_core_080 = input_i[0] & input_a[0];
  assign cgp_core_082 = ~(input_f[0] ^ input_h[1]);
  assign cgp_core_085 = input_e[1] | input_f[0];
  assign cgp_core_086 = ~(input_f[0] ^ input_a[1]);
  assign cgp_core_087 = cgp_core_082 | cgp_core_082;
  assign cgp_core_091 = ~input_g[1];
  assign cgp_core_095 = ~(input_e[1] ^ input_e[1]);
  assign cgp_core_096 = input_h[1] | input_b[1];
  assign cgp_core_099 = ~(input_b[0] & input_e[0]);
  assign cgp_core_101 = input_i[0] | cgp_core_096;
  assign cgp_core_104 = input_b[0] & input_d[1];
  assign cgp_core_105 = ~(input_e[1] & input_i[1]);
  assign cgp_core_107 = ~(input_i[1] & input_a[0]);

  assign cgp_out[0] = 1'b0;
endmodule