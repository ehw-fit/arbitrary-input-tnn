module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_032;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_072;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = input_d[1] ^ input_c[0];
  assign cgp_core_020 = input_d[0] | input_c[1];
  assign cgp_core_021 = ~input_a[2];
  assign cgp_core_026 = input_a[1] ^ input_c[2];
  assign cgp_core_027 = ~(input_b[0] & input_a[2]);
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_033_not = ~input_c[1];
  assign cgp_core_034 = ~(input_c[1] | input_e[2]);
  assign cgp_core_036 = input_d[2] ^ input_e[2];
  assign cgp_core_039 = input_b[1] & input_b[2];
  assign cgp_core_041 = ~(input_e[0] ^ input_d[0]);
  assign cgp_core_043 = input_e[0] ^ cgp_core_033_not;
  assign cgp_core_044 = cgp_core_021 & cgp_core_033_not;
  assign cgp_core_049 = input_a[1] & input_c[0];
  assign cgp_core_051 = input_c[1] & input_c[1];
  assign cgp_core_053 = ~(input_d[1] & input_e[1]);
  assign cgp_core_054 = ~(input_d[0] ^ input_c[2]);
  assign cgp_core_056 = cgp_core_053 & input_b[2];
  assign cgp_core_057 = cgp_core_054 | input_a[0];
  assign cgp_core_058 = ~(input_c[1] ^ input_d[0]);
  assign cgp_core_064 = input_a[0] & input_e[1];
  assign cgp_core_066 = ~input_c[0];
  assign cgp_core_068 = ~input_d[0];
  assign cgp_core_069 = input_c[1] & input_b[1];
  assign cgp_core_072 = input_e[1] & input_e[2];
  assign cgp_core_074_not = ~input_c[2];
  assign cgp_core_075 = ~(input_c[1] & cgp_core_072);
  assign cgp_core_076 = ~(input_d[2] ^ cgp_core_041);
  assign cgp_core_077 = ~(input_c[0] & input_a[2]);
  assign cgp_core_078 = ~(input_e[0] ^ input_b[1]);
  assign cgp_core_079 = input_c[1] | input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule