module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044_not;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080;

  assign cgp_core_019 = ~(input_a[2] ^ input_c[2]);
  assign cgp_core_020 = ~(input_c[2] ^ input_b[0]);
  assign cgp_core_021 = ~(input_b[2] ^ input_b[1]);
  assign cgp_core_023 = input_b[1] & input_b[1];
  assign cgp_core_024 = ~input_e[1];
  assign cgp_core_026_not = ~input_b[2];
  assign cgp_core_027 = input_b[1] & input_c[2];
  assign cgp_core_028 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_029 = ~(input_b[1] & input_a[2]);
  assign cgp_core_030 = input_a[0] | input_d[2];
  assign cgp_core_031 = input_d[0] & input_d[2];
  assign cgp_core_032 = input_a[2] & input_a[0];
  assign cgp_core_033 = ~(input_e[1] ^ input_e[1]);
  assign cgp_core_034 = input_a[1] | input_a[2];
  assign cgp_core_035 = ~input_b[2];
  assign cgp_core_037 = ~(input_a[1] ^ input_e[1]);
  assign cgp_core_038 = input_b[1] ^ input_a[2];
  assign cgp_core_039 = ~(input_a[0] ^ input_d[1]);
  assign cgp_core_040 = input_a[2] | input_a[2];
  assign cgp_core_041 = input_c[2] | input_b[2];
  assign cgp_core_042 = ~input_b[1];
  assign cgp_core_044_not = ~input_d[2];
  assign cgp_core_046 = ~(input_e[1] | input_b[0]);
  assign cgp_core_047 = ~(input_a[2] & input_d[0]);
  assign cgp_core_048 = input_c[1] | input_c[2];
  assign cgp_core_050 = ~input_d[2];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_055 = input_b[0] & input_c[1];
  assign cgp_core_056 = ~cgp_core_051;
  assign cgp_core_057 = cgp_core_041 & cgp_core_056;
  assign cgp_core_059 = ~(input_e[1] | input_b[2]);
  assign cgp_core_060 = input_a[1] | input_e[0];
  assign cgp_core_061 = ~input_d[1];
  assign cgp_core_062 = ~(input_a[1] | input_d[1]);
  assign cgp_core_063 = input_b[2] & input_c[2];
  assign cgp_core_064 = ~(input_e[1] ^ input_d[0]);
  assign cgp_core_065 = input_c[1] & input_e[1];
  assign cgp_core_067 = input_d[0] & input_c[1];
  assign cgp_core_071 = input_d[1] ^ input_d[2];
  assign cgp_core_073 = input_e[0] ^ input_a[2];
  assign cgp_core_076 = input_e[2] | cgp_core_063;
  assign cgp_core_077 = input_e[2] | cgp_core_076;
  assign cgp_core_078 = input_a[2] ^ input_e[1];
  assign cgp_core_080 = cgp_core_077 | cgp_core_057;

  assign cgp_out[0] = cgp_core_080;
endmodule