module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_071;

  assign cgp_core_014 = ~(input_f[0] | input_d[0]);
  assign cgp_core_015 = ~(input_c[1] & input_d[1]);
  assign cgp_core_016 = ~(input_d[1] & input_c[1]);
  assign cgp_core_019 = ~input_d[0];
  assign cgp_core_020 = ~(input_e[0] & input_b[0]);
  assign cgp_core_022_not = ~input_d[0];
  assign cgp_core_023 = ~(input_a[1] | input_d[1]);
  assign cgp_core_025_not = ~input_e[1];
  assign cgp_core_026 = ~(input_c[0] ^ input_e[1]);
  assign cgp_core_028 = ~input_c[0];
  assign cgp_core_029 = input_d[1] | input_d[1];
  assign cgp_core_032_not = ~input_e[1];
  assign cgp_core_033 = ~input_a[1];
  assign cgp_core_034_not = ~input_e[0];
  assign cgp_core_042 = ~input_c[0];
  assign cgp_core_045 = input_a[1] & input_e[1];
  assign cgp_core_054 = ~(input_a[0] ^ input_a[0]);
  assign cgp_core_055 = ~(input_a[1] | input_a[1]);
  assign cgp_core_056 = ~(input_d[1] ^ input_b[0]);
  assign cgp_core_057 = input_a[1] | input_c[0];
  assign cgp_core_062 = input_d[1] & input_e[1];
  assign cgp_core_063 = ~(input_e[1] ^ input_d[0]);
  assign cgp_core_064 = input_e[1] & input_e[1];
  assign cgp_core_065 = input_f[1] & input_e[0];
  assign cgp_core_066 = ~(input_b[0] & input_d[0]);
  assign cgp_core_067 = ~(input_b[1] | input_d[0]);
  assign cgp_core_069 = ~(input_c[0] & input_d[0]);
  assign cgp_core_071 = ~input_a[0];

  assign cgp_out[0] = 1'b1;
endmodule