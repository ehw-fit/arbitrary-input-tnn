module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_b[1] | input_c[0]);
  assign cgp_core_018 = ~(input_b[0] & input_d[0]);
  assign cgp_core_019 = ~input_e[0];
  assign cgp_core_024 = input_d[2] | input_d[2];
  assign cgp_core_026 = ~(input_c[0] & input_e[2]);
  assign cgp_core_027 = ~(input_a[1] ^ input_b[1]);
  assign cgp_core_028 = input_c[1] | input_a[1];
  assign cgp_core_029 = ~input_c[0];
  assign cgp_core_031 = input_e[2] | input_a[2];
  assign cgp_core_032 = input_d[1] & input_b[0];
  assign cgp_core_033 = input_b[0] | input_d[1];
  assign cgp_core_035 = ~input_a[1];
  assign cgp_core_036 = ~input_b[2];
  assign cgp_core_037 = input_d[2] ^ input_b[0];
  assign cgp_core_039 = input_d[1] ^ input_b[2];
  assign cgp_core_041 = ~input_d[2];
  assign cgp_core_045 = input_a[0] ^ input_c[2];
  assign cgp_core_048 = input_c[0] ^ input_b[1];
  assign cgp_core_049 = ~(cgp_core_026 & input_e[2]);
  assign cgp_core_050 = ~(input_e[2] | input_c[0]);
  assign cgp_core_051 = input_c[2] & input_b[1];
  assign cgp_core_055 = input_a[1] ^ input_d[1];
  assign cgp_core_057 = input_e[0] | input_a[0];
  assign cgp_core_058 = ~(input_a[2] & input_c[0]);
  assign cgp_core_059 = ~(input_d[2] & input_c[1]);
  assign cgp_core_061 = cgp_core_055 & input_e[0];
  assign cgp_core_062 = cgp_core_061 & input_d[2];
  assign cgp_core_063 = input_a[0] | input_c[1];
  assign cgp_core_064 = input_a[1] | input_a[2];
  assign cgp_core_066 = ~input_d[0];
  assign cgp_core_068 = ~(input_c[2] & cgp_core_045);
  assign cgp_core_069 = input_e[1] ^ input_b[1];
  assign cgp_core_070 = input_e[1] & input_d[2];
  assign cgp_core_072 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_073 = ~(input_d[1] ^ input_d[0]);
  assign cgp_core_075 = ~(input_e[0] & cgp_core_072);
  assign cgp_core_076 = ~input_c[1];
  assign cgp_core_079 = input_c[1] ^ input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule