module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_052_not;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_089;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_097;
  wire cgp_core_098;

  assign cgp_core_024 = input_c[1] ^ input_b[1];
  assign cgp_core_026 = input_f[1] ^ input_e[1];
  assign cgp_core_027 = ~(input_c[0] ^ input_c[0]);
  assign cgp_core_029 = ~(input_a[0] | input_e[2]);
  assign cgp_core_030 = ~input_b[2];
  assign cgp_core_032 = ~(input_d[1] & input_a[1]);
  assign cgp_core_033 = ~(input_b[0] | input_d[1]);
  assign cgp_core_034 = input_e[1] & input_c[2];
  assign cgp_core_035 = ~(input_b[0] & input_a[2]);
  assign cgp_core_036 = ~(input_e[0] ^ input_d[0]);
  assign cgp_core_037 = ~(input_e[2] | input_b[2]);
  assign cgp_core_038 = ~(input_c[1] | input_d[1]);
  assign cgp_core_042 = ~input_c[0];
  assign cgp_core_043 = input_a[2] ^ input_b[0];
  assign cgp_core_044 = input_c[0] & input_a[1];
  assign cgp_core_045 = ~(input_d[0] | input_e[1]);
  assign cgp_core_047 = ~input_d[2];
  assign cgp_core_052_not = ~input_a[1];
  assign cgp_core_054 = ~input_d[1];
  assign cgp_core_056 = input_d[1] & input_f[0];
  assign cgp_core_057 = ~(input_a[1] & input_f[0]);
  assign cgp_core_059 = ~(input_c[0] & input_a[2]);
  assign cgp_core_060 = input_e[0] ^ input_c[1];
  assign cgp_core_063 = input_b[2] & input_b[0];
  assign cgp_core_064 = ~(input_a[0] ^ input_f[1]);
  assign cgp_core_070 = input_b[0] | input_f[2];
  assign cgp_core_071 = input_a[2] | input_b[0];
  assign cgp_core_074 = input_c[2] & input_f[2];
  assign cgp_core_075 = ~(input_c[0] | input_e[0]);
  assign cgp_core_077 = input_a[2] & input_c[2];
  assign cgp_core_080 = ~(input_b[1] | input_d[1]);
  assign cgp_core_081 = ~(input_b[1] | input_d[2]);
  assign cgp_core_082 = input_b[2] ^ input_c[0];
  assign cgp_core_083 = ~(input_b[1] ^ input_a[1]);
  assign cgp_core_085 = ~(input_d[2] & input_d[0]);
  assign cgp_core_086 = ~input_e[2];
  assign cgp_core_089 = input_a[0] | input_f[2];
  assign cgp_core_093 = ~input_e[0];
  assign cgp_core_094 = ~(input_b[1] & input_b[1]);
  assign cgp_core_097 = ~(input_e[2] | input_d[0]);
  assign cgp_core_098 = cgp_core_077 | input_e[2];

  assign cgp_out[0] = cgp_core_098;
endmodule