module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_034_not;
  wire cgp_core_037_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060_not;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_016 = input_g[1] & input_e[0];
  assign cgp_core_017 = ~(input_c[0] ^ input_a[0]);
  assign cgp_core_018 = input_a[0] | input_b[0];
  assign cgp_core_019 = input_b[1] ^ input_c[0];
  assign cgp_core_020 = ~(input_e[1] & input_b[1]);
  assign cgp_core_021 = input_f[0] ^ input_f[0];
  assign cgp_core_023 = ~(input_a[1] & input_c[0]);
  assign cgp_core_024 = input_f[0] ^ input_b[0];
  assign cgp_core_026 = ~(input_a[1] | input_d[1]);
  assign cgp_core_029 = ~(input_c[1] | input_a[0]);
  assign cgp_core_031 = input_e[1] & input_a[1];
  assign cgp_core_034_not = ~input_d[0];
  assign cgp_core_037_not = ~input_a[1];
  assign cgp_core_038 = input_a[1] & input_f[0];
  assign cgp_core_039 = ~input_b[1];
  assign cgp_core_040 = ~(input_b[1] & input_e[1]);
  assign cgp_core_042 = input_a[1] ^ input_b[1];
  assign cgp_core_043 = input_b[1] | input_c[1];
  assign cgp_core_045 = ~(input_e[1] & input_e[0]);
  assign cgp_core_046 = ~(input_a[0] ^ input_f[0]);
  assign cgp_core_048 = ~(input_e[1] | input_b[1]);
  assign cgp_core_049 = input_c[0] ^ input_d[1];
  assign cgp_core_050_not = ~input_c[1];
  assign cgp_core_051 = ~(input_c[1] ^ input_e[1]);
  assign cgp_core_054 = input_a[1] | input_g[0];
  assign cgp_core_055 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_057 = input_d[1] | input_g[0];
  assign cgp_core_058 = input_c[1] & input_a[0];
  assign cgp_core_059 = cgp_core_031 & input_d[1];
  assign cgp_core_060_not = ~input_b[1];
  assign cgp_core_061 = input_e[1] ^ input_f[1];
  assign cgp_core_062 = ~(input_e[1] | input_a[1]);
  assign cgp_core_063 = ~(input_f[0] | input_f[0]);
  assign cgp_core_064 = input_a[1] & input_d[1];
  assign cgp_core_065 = ~input_b[1];
  assign cgp_core_066 = ~(input_f[1] ^ input_d[1]);
  assign cgp_core_067 = ~(input_f[1] | input_d[0]);
  assign cgp_core_068 = ~(input_b[0] | input_a[0]);
  assign cgp_core_069 = ~(input_c[1] | input_e[0]);
  assign cgp_core_070 = ~input_b[1];
  assign cgp_core_072 = ~input_g[0];
  assign cgp_core_073 = ~(input_a[1] & input_g[1]);
  assign cgp_core_075 = input_f[0] ^ input_f[0];
  assign cgp_core_076 = ~input_e[1];
  assign cgp_core_077 = ~(input_f[0] | input_f[1]);
  assign cgp_core_079 = ~(input_e[1] | input_e[0]);

  assign cgp_out[0] = cgp_core_059;
endmodule