module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = ~(input_f[0] | input_e[0]);
  assign cgp_core_017 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_018 = input_b[1] | input_a[1];
  assign cgp_core_019 = ~(input_c[1] ^ input_b[1]);
  assign cgp_core_020 = input_d[0] ^ input_b[1];
  assign cgp_core_021 = ~input_b[1];
  assign cgp_core_023 = ~(input_e[0] & input_f[1]);
  assign cgp_core_024 = ~(input_a[0] ^ input_f[1]);
  assign cgp_core_025 = ~(input_d[0] ^ input_a[1]);
  assign cgp_core_027 = ~(input_c[0] & input_f[0]);
  assign cgp_core_031 = input_a[1] & input_d[1];
  assign cgp_core_032 = ~input_g[1];
  assign cgp_core_036 = ~(input_f[1] | input_g[0]);
  assign cgp_core_037 = input_g[0] & input_b[1];
  assign cgp_core_038 = input_b[0] & input_f[0];
  assign cgp_core_039 = ~(input_e[0] ^ input_b[1]);
  assign cgp_core_041 = ~(input_e[1] ^ input_c[1]);
  assign cgp_core_043 = ~input_d[1];
  assign cgp_core_044 = ~(input_a[0] | input_g[0]);
  assign cgp_core_046_not = ~input_f[0];
  assign cgp_core_049 = ~(input_a[0] | input_a[1]);
  assign cgp_core_050 = ~(input_g[0] & input_g[1]);
  assign cgp_core_053 = input_e[1] & input_c[1];
  assign cgp_core_054 = cgp_core_038 & input_g[1];
  assign cgp_core_055_not = ~input_b[1];
  assign cgp_core_056 = input_c[1] & input_f[1];
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = cgp_core_031 & cgp_core_058;
  assign cgp_core_060 = ~(input_b[1] | cgp_core_057);
  assign cgp_core_061 = ~(input_b[0] | input_b[0]);
  assign cgp_core_062 = ~(input_g[1] | input_b[0]);
  assign cgp_core_063 = input_e[1] & cgp_core_060;
  assign cgp_core_064 = input_a[1] | input_a[0];
  assign cgp_core_065 = input_e[0] | input_c[1];
  assign cgp_core_069 = input_f[1] | input_a[1];
  assign cgp_core_070 = input_c[0] & input_b[0];
  assign cgp_core_071 = ~(input_f[1] | input_f[1]);
  assign cgp_core_072 = input_c[0] ^ input_b[1];
  assign cgp_core_074 = ~input_b[0];
  assign cgp_core_076 = ~input_e[1];
  assign cgp_core_078 = cgp_core_063 | cgp_core_059;
  assign cgp_core_079 = ~(input_f[1] & input_f[1]);

  assign cgp_out[0] = cgp_core_078;
endmodule