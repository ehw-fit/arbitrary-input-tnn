module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012_not;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031_not;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_054;

  assign cgp_core_012_not = ~input_e[1];
  assign cgp_core_013 = input_d[0] & input_b[0];
  assign cgp_core_014 = input_b[1] | input_d[1];
  assign cgp_core_015 = input_b[1] & input_d[1];
  assign cgp_core_017 = cgp_core_014 & cgp_core_013;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~(input_a[1] ^ input_b[1]);
  assign cgp_core_020 = ~input_b[1];
  assign cgp_core_021 = input_c[1] | input_e[1];
  assign cgp_core_022 = input_c[1] & input_e[1];
  assign cgp_core_024 = input_d[1] | input_b[1];
  assign cgp_core_026 = input_c[0] ^ input_a[0];
  assign cgp_core_029 = input_a[1] & cgp_core_021;
  assign cgp_core_030 = ~(input_e[0] ^ input_e[1]);
  assign cgp_core_031_not = ~input_b[0];
  assign cgp_core_033 = cgp_core_022 | cgp_core_029;
  assign cgp_core_034_not = ~input_c[1];
  assign cgp_core_037 = ~cgp_core_033;
  assign cgp_core_038 = cgp_core_018 & cgp_core_037;
  assign cgp_core_040 = ~(input_c[1] | input_a[1]);
  assign cgp_core_042 = ~input_e[1];
  assign cgp_core_043 = cgp_core_014 & cgp_core_042;
  assign cgp_core_044 = cgp_core_043 & cgp_core_040;
  assign cgp_core_046 = input_a[1] | input_e[1];
  assign cgp_core_047 = ~(input_c[0] & input_d[0]);
  assign cgp_core_049 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_050 = input_e[0] ^ input_a[1];
  assign cgp_core_051 = ~(input_b[0] | input_d[0]);
  assign cgp_core_054 = cgp_core_044 | cgp_core_038;

  assign cgp_out[0] = cgp_core_054;
endmodule