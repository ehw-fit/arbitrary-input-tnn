module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058_not;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062_not;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086_not;
  wire cgp_core_087;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;

  assign cgp_core_019 = input_d[0] & input_c[1];
  assign cgp_core_020 = ~(input_h[1] | input_h[0]);
  assign cgp_core_021 = input_e[0] & input_b[1];
  assign cgp_core_022 = ~input_f[1];
  assign cgp_core_023_not = ~input_c[1];
  assign cgp_core_024 = input_h[0] | input_h[1];
  assign cgp_core_025 = ~(input_b[1] ^ input_g[0]);
  assign cgp_core_026 = ~(input_b[0] & input_d[0]);
  assign cgp_core_027 = ~input_h[0];
  assign cgp_core_028 = ~(input_a[1] ^ input_g[1]);
  assign cgp_core_031 = input_a[0] ^ input_c[0];
  assign cgp_core_034 = input_b[1] | input_e[1];
  assign cgp_core_035 = ~(input_b[0] | input_h[1]);
  assign cgp_core_036 = input_c[1] | input_b[1];
  assign cgp_core_037 = ~(input_h[0] ^ input_c[0]);
  assign cgp_core_038 = input_c[1] ^ input_f[0];
  assign cgp_core_040 = ~(input_f[1] | input_b[0]);
  assign cgp_core_041 = input_f[0] | input_c[1];
  assign cgp_core_043 = input_e[0] ^ input_h[1];
  assign cgp_core_045 = input_g[1] ^ input_d[1];
  assign cgp_core_049 = input_c[0] ^ input_g[1];
  assign cgp_core_051 = ~(input_a[1] | input_c[0]);
  assign cgp_core_052 = input_e[1] ^ input_a[1];
  assign cgp_core_053 = ~(input_f[0] | input_e[1]);
  assign cgp_core_054 = ~(input_b[1] | input_e[0]);
  assign cgp_core_055 = input_c[0] & input_e[0];
  assign cgp_core_057 = ~(input_g[1] | input_f[0]);
  assign cgp_core_058_not = ~input_b[0];
  assign cgp_core_060 = ~(input_b[0] & input_a[1]);
  assign cgp_core_061 = ~input_g[0];
  assign cgp_core_062_not = ~input_h[0];
  assign cgp_core_063 = ~(input_e[1] | input_b[1]);
  assign cgp_core_064 = ~input_d[0];
  assign cgp_core_065 = input_b[1] & input_g[0];
  assign cgp_core_066 = ~input_h[0];
  assign cgp_core_067 = ~(input_h[0] | input_g[0]);
  assign cgp_core_068 = ~(input_e[0] & input_f[1]);
  assign cgp_core_069 = ~(input_c[0] ^ input_a[1]);
  assign cgp_core_078 = input_c[0] & input_c[0];
  assign cgp_core_079 = ~(input_c[1] & input_d[0]);
  assign cgp_core_080 = input_f[1] | input_f[0];
  assign cgp_core_081 = ~(input_b[1] & input_d[0]);
  assign cgp_core_082 = input_c[1] & input_e[0];
  assign cgp_core_083 = ~(input_f[1] ^ input_b[1]);
  assign cgp_core_085 = ~(input_f[0] ^ input_b[1]);
  assign cgp_core_086_not = ~input_f[1];
  assign cgp_core_087 = input_f[1] | input_a[1];
  assign cgp_core_091 = ~(input_b[0] ^ input_g[1]);
  assign cgp_core_092 = ~(input_f[1] | input_a[0]);
  assign cgp_core_093 = input_a[1] | input_b[0];
  assign cgp_core_094 = ~(input_c[1] ^ input_a[0]);

  assign cgp_out[0] = 1'b0;
endmodule