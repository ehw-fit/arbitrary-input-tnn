module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047_not;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078_not;
  wire cgp_core_080;
  wire cgp_core_083;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089_not;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;
  wire cgp_core_095;

  assign cgp_core_022 = input_a[1] & input_b[1];
  assign cgp_core_023 = input_b[1] & input_b[1];
  assign cgp_core_024 = ~(input_b[0] | input_c[2]);
  assign cgp_core_025 = input_e[1] | input_b[0];
  assign cgp_core_026 = ~(input_f[1] | input_c[1]);
  assign cgp_core_027 = ~(input_a[1] ^ input_f[0]);
  assign cgp_core_028 = input_f[2] | input_c[1];
  assign cgp_core_029 = ~(cgp_core_027 ^ cgp_core_026);
  assign cgp_core_030 = input_f[1] | cgp_core_026;
  assign cgp_core_031 = ~input_f[0];
  assign cgp_core_034 = input_c[1] | input_d[1];
  assign cgp_core_035 = input_d[2] ^ input_c[2];
  assign cgp_core_037 = ~cgp_core_034;
  assign cgp_core_038 = input_a[1] | input_b[1];
  assign cgp_core_039 = input_b[2] ^ input_d[2];
  assign cgp_core_041 = ~cgp_core_039;
  assign cgp_core_042 = input_c[2] & cgp_core_038;
  assign cgp_core_043 = input_f[1] | input_e[0];
  assign cgp_core_045 = ~(input_a[1] & input_f[0]);
  assign cgp_core_046 = ~(input_d[0] & input_e[0]);
  assign cgp_core_047_not = ~input_f[1];
  assign cgp_core_048 = ~(input_f[1] ^ input_a[1]);
  assign cgp_core_050 = ~(input_e[0] & input_f[0]);
  assign cgp_core_053 = input_d[1] & input_b[0];
  assign cgp_core_055 = ~(input_c[2] & input_e[0]);
  assign cgp_core_057 = input_a[2] & input_f[2];
  assign cgp_core_058 = input_a[1] ^ input_a[1];
  assign cgp_core_060 = input_a[0] & input_e[0];
  assign cgp_core_061 = ~(input_c[0] & input_b[1]);
  assign cgp_core_062 = input_b[0] | input_f[2];
  assign cgp_core_063 = input_d[2] ^ input_c[0];
  assign cgp_core_065 = ~(input_c[1] ^ cgp_core_062);
  assign cgp_core_066 = ~(input_d[1] ^ input_b[1]);
  assign cgp_core_067 = ~(input_f[2] ^ input_f[1]);
  assign cgp_core_068 = input_c[0] ^ cgp_core_055;
  assign cgp_core_069 = input_b[1] | cgp_core_055;
  assign cgp_core_071 = input_c[0] | input_c[1];
  assign cgp_core_075 = ~input_f[0];
  assign cgp_core_077 = input_e[0] & input_e[2];
  assign cgp_core_078_not = ~input_f[2];
  assign cgp_core_080 = input_b[2] ^ cgp_core_065;
  assign cgp_core_083 = input_e[1] | cgp_core_065;
  assign cgp_core_086 = cgp_core_024 ^ input_e[1];
  assign cgp_core_088 = cgp_core_024 ^ input_e[0];
  assign cgp_core_089_not = ~input_a[0];
  assign cgp_core_090 = ~input_a[0];
  assign cgp_core_091 = input_e[1] & cgp_core_090;
  assign cgp_core_093 = ~(input_b[0] | input_a[2]);
  assign cgp_core_095 = ~(input_a[0] | input_f[0]);

  assign cgp_out[0] = 1'b0;
endmodule