module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058_not;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_088;

  assign cgp_core_023 = input_a[1] & input_d[2];
  assign cgp_core_027 = ~input_a[0];
  assign cgp_core_028 = input_a[2] & input_d[1];
  assign cgp_core_030 = ~cgp_core_027;
  assign cgp_core_031 = input_a[1] | cgp_core_030;
  assign cgp_core_032 = ~input_c[0];
  assign cgp_core_033 = input_c[0] & input_d[0];
  assign cgp_core_035 = ~input_c[1];
  assign cgp_core_036_not = ~cgp_core_033;
  assign cgp_core_038 = input_c[0] | input_f[0];
  assign cgp_core_039 = input_c[2] ^ input_d[2];
  assign cgp_core_040 = input_c[2] & input_b[2];
  assign cgp_core_041 = ~(cgp_core_039 | input_a[1]);
  assign cgp_core_042 = cgp_core_039 & input_c[2];
  assign cgp_core_043 = ~(input_a[1] | input_e[0]);
  assign cgp_core_046 = input_e[1] ^ input_f[1];
  assign cgp_core_047 = input_e[1] & input_f[1];
  assign cgp_core_048 = cgp_core_046 ^ input_e[0];
  assign cgp_core_049 = cgp_core_046 & input_e[0];
  assign cgp_core_050 = cgp_core_047 | cgp_core_049;
  assign cgp_core_051 = input_e[2] ^ input_f[2];
  assign cgp_core_052 = input_e[2] & input_f[2];
  assign cgp_core_053 = cgp_core_051 ^ cgp_core_050;
  assign cgp_core_054 = ~input_b[1];
  assign cgp_core_055 = cgp_core_052 | cgp_core_054;
  assign cgp_core_057 = cgp_core_032 & input_e[0];
  assign cgp_core_058_not = ~cgp_core_048;
  assign cgp_core_059 = cgp_core_036_not & cgp_core_048;
  assign cgp_core_061 = ~cgp_core_058_not;
  assign cgp_core_062 = input_b[2] | cgp_core_061;
  assign cgp_core_063 = cgp_core_041 ^ cgp_core_053;
  assign cgp_core_064 = cgp_core_041 & cgp_core_053;
  assign cgp_core_065 = input_f[2] ^ cgp_core_062;
  assign cgp_core_068 = cgp_core_043 | input_d[1];
  assign cgp_core_069 = input_b[0] & input_f[2];
  assign cgp_core_070 = cgp_core_068 ^ input_f[1];
  assign cgp_core_072 = input_a[0] | cgp_core_068;
  assign cgp_core_073 = ~(cgp_core_072 & cgp_core_072);
  assign cgp_core_074 = ~cgp_core_072;
  assign cgp_core_075 = input_d[2] ^ cgp_core_070;
  assign cgp_core_078 = ~(input_b[0] ^ cgp_core_070);
  assign cgp_core_080 = ~cgp_core_065;
  assign cgp_core_088 = ~(input_a[0] | input_d[2]);

  assign cgp_out[0] = 1'b0;
endmodule