module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_014 = input_a[0] ^ input_c[0];
  assign cgp_core_016 = ~(input_a[0] & input_e[0]);
  assign cgp_core_020 = input_f[0] & input_c[0];
  assign cgp_core_021 = ~input_e[1];
  assign cgp_core_022 = input_d[1] & input_c[0];
  assign cgp_core_024_not = ~input_f[0];
  assign cgp_core_025 = input_d[0] | input_a[0];
  assign cgp_core_028 = input_a[0] & input_d[0];
  assign cgp_core_029_not = ~input_f[1];
  assign cgp_core_030 = ~(input_e[1] ^ input_b[1]);
  assign cgp_core_031 = ~(input_d[0] | input_c[0]);
  assign cgp_core_033 = ~input_b[1];
  assign cgp_core_034 = ~input_d[1];
  assign cgp_core_036 = input_d[0] & input_f[0];
  assign cgp_core_037 = ~cgp_core_014;
  assign cgp_core_039 = input_a[0] | input_d[1];
  assign cgp_core_040 = input_a[0] & input_d[1];
  assign cgp_core_041 = cgp_core_039 | input_c[0];
  assign cgp_core_042 = input_d[1] & input_c[0];
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;
  assign cgp_core_044 = input_a[1] | input_e[0];
  assign cgp_core_045 = ~input_d[0];
  assign cgp_core_046 = cgp_core_044 | cgp_core_043;
  assign cgp_core_048 = input_d[0] & input_e[0];
  assign cgp_core_049 = cgp_core_036 | input_f[1];
  assign cgp_core_050 = ~(input_e[1] & input_b[0]);
  assign cgp_core_053 = ~(input_b[1] ^ input_a[1]);
  assign cgp_core_054 = input_c[1] & input_d[0];
  assign cgp_core_056 = ~input_b[0];
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_059 = cgp_core_041 & cgp_core_058;
  assign cgp_core_061 = ~(cgp_core_041 ^ input_b[1]);
  assign cgp_core_062 = cgp_core_061 & cgp_core_056;
  assign cgp_core_065 = input_e[1] | input_f[0];
  assign cgp_core_067 = cgp_core_037 & cgp_core_062;
  assign cgp_core_068 = cgp_core_059 | cgp_core_046;
  assign cgp_core_069 = input_c[1] | cgp_core_068;
  assign cgp_core_070 = input_e[1] | cgp_core_067;
  assign cgp_core_071 = cgp_core_049 | cgp_core_070;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;

  assign cgp_out[0] = cgp_core_072;
endmodule