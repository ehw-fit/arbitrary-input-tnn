module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;

  assign cgp_core_018 = input_b[0] | input_h[0];
  assign cgp_core_019 = ~(input_d[0] | input_g[1]);
  assign cgp_core_020 = ~input_h[1];
  assign cgp_core_021 = input_d[1] & input_h[1];
  assign cgp_core_022 = input_a[0] ^ input_h[1];
  assign cgp_core_023 = cgp_core_020 & input_g[0];
  assign cgp_core_025 = ~input_h[1];
  assign cgp_core_027 = input_d[0] ^ input_c[1];
  assign cgp_core_028_not = ~input_h[1];
  assign cgp_core_029 = input_g[0] ^ input_c[0];
  assign cgp_core_032 = ~input_c[1];
  assign cgp_core_034 = input_b[0] ^ input_a[0];
  assign cgp_core_035 = input_b[0] | input_d[0];
  assign cgp_core_036 = ~(input_e[0] | input_f[1]);
  assign cgp_core_037 = input_b[1] & input_c[1];
  assign cgp_core_038 = input_c[0] ^ input_e[1];
  assign cgp_core_039 = cgp_core_036 & cgp_core_035;
  assign cgp_core_040 = input_f[0] | input_a[0];
  assign cgp_core_041 = input_f[0] ^ input_d[1];
  assign cgp_core_044 = input_b[1] & input_h[1];
  assign cgp_core_047 = ~cgp_core_044;
  assign cgp_core_048 = input_e[0] ^ cgp_core_041;
  assign cgp_core_049 = ~(input_d[1] & cgp_core_041);
  assign cgp_core_052 = ~input_f[0];
  assign cgp_core_053 = input_f[0] ^ input_d[0];
  assign cgp_core_054 = ~(input_h[1] | input_f[1]);
  assign cgp_core_055 = cgp_core_047 & input_e[0];
  assign cgp_core_058 = cgp_core_034 & cgp_core_048;
  assign cgp_core_059 = ~(cgp_core_038 ^ input_c[0]);
  assign cgp_core_060 = cgp_core_038 & cgp_core_052;
  assign cgp_core_061 = cgp_core_059 ^ cgp_core_058;
  assign cgp_core_062 = input_a[1] & input_b[0];
  assign cgp_core_065 = input_f[0] & cgp_core_055;
  assign cgp_core_066 = input_c[1] & input_e[0];
  assign cgp_core_067 = ~input_g[0];
  assign cgp_core_069 = input_g[1] ^ input_b[1];
  assign cgp_core_071 = ~input_b[0];
  assign cgp_core_072 = ~input_a[1];
  assign cgp_core_073 = input_b[0] ^ input_g[1];
  assign cgp_core_078 = ~(input_f[0] | cgp_core_066);
  assign cgp_core_079 = ~(input_b[0] & cgp_core_078);
  assign cgp_core_083 = ~cgp_core_061;
  assign cgp_core_084 = cgp_core_029 ^ cgp_core_083;
  assign cgp_core_085 = input_d[0] & input_b[1];
  assign cgp_core_088 = ~input_c[0];
  assign cgp_core_089 = ~input_c[0];
  assign cgp_core_090 = input_e[0] & input_c[0];

  assign cgp_out[0] = 1'b0;
endmodule