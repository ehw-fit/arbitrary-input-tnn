module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_033_not;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;

  assign cgp_core_014 = input_a[5] & input_a[8];
  assign cgp_core_015 = ~(input_a[4] & input_a[2]);
  assign cgp_core_016 = input_a[8] ^ input_a[9];
  assign cgp_core_017 = ~input_a[3];
  assign cgp_core_019 = ~(input_a[7] & input_a[11]);
  assign cgp_core_020 = ~(input_a[7] | input_a[1]);
  assign cgp_core_023 = input_a[10] | input_a[3];
  assign cgp_core_024 = input_a[4] ^ input_a[6];
  assign cgp_core_025 = ~input_a[4];
  assign cgp_core_026 = ~(input_a[6] & input_a[4]);
  assign cgp_core_027 = input_a[2] & input_a[1];
  assign cgp_core_029 = ~(input_a[3] ^ input_a[2]);
  assign cgp_core_033_not = ~input_a[10];
  assign cgp_core_035 = ~(input_a[5] | input_a[2]);
  assign cgp_core_036 = input_a[4] | input_a[3];
  assign cgp_core_038 = input_a[2] ^ input_a[7];
  assign cgp_core_040 = input_a[5] & input_a[3];
  assign cgp_core_042 = ~(input_a[6] & input_a[3]);
  assign cgp_core_043 = input_a[0] | input_a[4];
  assign cgp_core_044 = ~(input_a[3] ^ input_a[5]);
  assign cgp_core_047 = input_a[5] | input_a[11];
  assign cgp_core_048 = input_a[9] ^ input_a[11];
  assign cgp_core_051 = input_a[9] | input_a[7];
  assign cgp_core_052 = ~(input_a[5] & input_a[10]);
  assign cgp_core_053 = input_a[10] | input_a[5];
  assign cgp_core_055_not = ~input_a[10];
  assign cgp_core_056 = ~(input_a[1] | input_a[5]);
  assign cgp_core_057 = ~(input_a[1] | input_a[9]);
  assign cgp_core_059 = ~input_a[11];
  assign cgp_core_060 = input_a[2] & input_a[8];
  assign cgp_core_061 = input_a[4] ^ input_a[8];
  assign cgp_core_063 = input_a[4] ^ input_a[5];
  assign cgp_core_064 = input_a[7] ^ input_a[10];
  assign cgp_core_070 = ~input_a[6];
  assign cgp_core_071 = input_a[7] & input_a[7];
  assign cgp_core_073 = ~(input_a[0] | input_a[7]);
  assign cgp_core_074 = ~(input_a[10] | input_a[3]);
  assign cgp_core_075 = input_a[11] | input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[3];
  assign cgp_core_077 = input_a[8] ^ input_a[9];

  assign cgp_out[0] = 1'b1;
  assign cgp_out[1] = 1'b1;
  assign cgp_out[2] = input_a[0];
  assign cgp_out[3] = 1'b0;
endmodule