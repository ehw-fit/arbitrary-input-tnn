module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_102;
  wire cgp_core_105_not;
  wire cgp_core_106;
  wire cgp_core_110;

  assign cgp_core_020 = input_c[0] & input_b[1];
  assign cgp_core_023_not = ~input_e[1];
  assign cgp_core_024 = ~(input_c[0] & input_a[0]);
  assign cgp_core_027 = ~(input_e[1] | input_i[1]);
  assign cgp_core_029 = input_g[1] ^ input_h[0];
  assign cgp_core_030 = ~(input_b[0] | input_h[1]);
  assign cgp_core_034 = ~(input_f[1] | input_f[0]);
  assign cgp_core_035 = input_i[1] & input_d[1];
  assign cgp_core_039 = ~(input_a[0] ^ input_e[1]);
  assign cgp_core_040 = input_e[1] & input_g[1];
  assign cgp_core_046 = input_i[0] & input_e[0];
  assign cgp_core_047 = input_g[0] | input_d[1];
  assign cgp_core_048 = ~input_c[1];
  assign cgp_core_049 = ~(input_b[0] ^ input_f[0]);
  assign cgp_core_050 = input_f[1] | input_a[1];
  assign cgp_core_055 = ~(input_d[1] | input_e[1]);
  assign cgp_core_056 = ~(input_i[1] ^ input_a[1]);
  assign cgp_core_061 = ~(input_e[1] & input_h[0]);
  assign cgp_core_062 = input_f[1] | input_a[1];
  assign cgp_core_063 = input_g[1] | input_e[0];
  assign cgp_core_064 = input_g[1] | input_i[1];
  assign cgp_core_065 = input_c[0] ^ input_b[0];
  assign cgp_core_066 = input_g[1] | input_b[1];
  assign cgp_core_067 = ~(input_h[1] ^ input_e[1]);
  assign cgp_core_068 = ~(input_e[0] ^ input_e[1]);
  assign cgp_core_069 = ~(input_e[1] | input_d[1]);
  assign cgp_core_071 = input_h[1] | input_d[1];
  assign cgp_core_072 = ~input_e[0];
  assign cgp_core_075 = cgp_core_050 ^ cgp_core_066;
  assign cgp_core_076 = ~(input_g[0] & input_h[1]);
  assign cgp_core_077 = ~cgp_core_075;
  assign cgp_core_079 = input_b[1] | cgp_core_075;
  assign cgp_core_081 = input_h[1] ^ input_c[1];
  assign cgp_core_082 = input_g[1] | cgp_core_079;
  assign cgp_core_083 = input_c[0] & input_e[1];
  assign cgp_core_084 = input_g[0] ^ input_d[1];
  assign cgp_core_085 = input_b[0] | input_e[0];
  assign cgp_core_086 = input_f[0] | input_e[0];
  assign cgp_core_087 = ~cgp_core_082;
  assign cgp_core_088 = cgp_core_035 & cgp_core_087;
  assign cgp_core_094 = ~(input_i[1] ^ input_f[0]);
  assign cgp_core_095 = ~(input_c[1] | cgp_core_077);
  assign cgp_core_096 = cgp_core_095 & cgp_core_035;
  assign cgp_core_097 = input_h[0] ^ input_h[0];
  assign cgp_core_099 = input_h[1] & cgp_core_096;
  assign cgp_core_100 = input_i[1] | input_i[1];
  assign cgp_core_102 = input_g[0] | input_c[1];
  assign cgp_core_105_not = ~input_g[0];
  assign cgp_core_106 = ~(input_h[1] ^ input_e[1]);
  assign cgp_core_110 = cgp_core_099 | cgp_core_088;

  assign cgp_out[0] = cgp_core_110;
endmodule