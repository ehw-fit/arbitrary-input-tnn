module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_020_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051_not;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068_not;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;

  assign cgp_core_016 = input_c[0] ^ input_e[1];
  assign cgp_core_020_not = ~input_d[0];
  assign cgp_core_024 = input_e[0] & input_g[0];
  assign cgp_core_025 = ~input_e[1];
  assign cgp_core_028 = ~(cgp_core_025 & cgp_core_024);
  assign cgp_core_029 = input_d[1] | input_e[0];
  assign cgp_core_031 = ~(cgp_core_016 & input_b[0]);
  assign cgp_core_032 = cgp_core_020_not ^ input_f[1];
  assign cgp_core_033 = input_a[1] & input_b[0];
  assign cgp_core_034 = cgp_core_032 ^ input_e[1];
  assign cgp_core_035_not = ~cgp_core_031;
  assign cgp_core_036 = cgp_core_033 | cgp_core_035_not;
  assign cgp_core_038 = ~(input_b[1] & cgp_core_029);
  assign cgp_core_039 = ~(cgp_core_029 | cgp_core_036);
  assign cgp_core_040 = ~cgp_core_029;
  assign cgp_core_042 = ~(input_b[0] ^ input_f[0]);
  assign cgp_core_043 = ~(input_g[0] ^ input_f[0]);
  assign cgp_core_044 = ~input_b[1];
  assign cgp_core_046 = input_c[0] ^ cgp_core_043;
  assign cgp_core_048 = ~(input_a[1] & input_d[1]);
  assign cgp_core_049 = input_f[1] ^ cgp_core_042;
  assign cgp_core_050 = input_a[0] & cgp_core_042;
  assign cgp_core_051_not = ~cgp_core_046;
  assign cgp_core_052 = input_c[1] & cgp_core_046;
  assign cgp_core_055 = cgp_core_052 | input_c[1];
  assign cgp_core_056 = ~(input_g[1] ^ input_a[1]);
  assign cgp_core_057 = ~(cgp_core_048 | cgp_core_055);
  assign cgp_core_058 = ~(cgp_core_057 & input_f[1]);
  assign cgp_core_061 = ~cgp_core_056;
  assign cgp_core_062 = cgp_core_039 & cgp_core_061;
  assign cgp_core_064 = ~(cgp_core_039 ^ cgp_core_056);
  assign cgp_core_067 = ~input_f[0];
  assign cgp_core_068_not = ~input_c[0];
  assign cgp_core_069_not = ~cgp_core_034;
  assign cgp_core_070 = input_d[0] & input_e[1];
  assign cgp_core_073 = input_d[1] & input_f[0];
  assign cgp_core_076 = cgp_core_073 & input_c[0];
  assign cgp_core_077 = input_e[1] | cgp_core_070;

  assign cgp_out[0] = 1'b1;
endmodule