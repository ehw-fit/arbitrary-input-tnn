module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_088;
  wire cgp_core_089;

  assign cgp_core_016 = input_a[12] ^ input_a[5];
  assign cgp_core_017 = ~(input_a[4] | input_a[0]);
  assign cgp_core_020 = ~(input_a[9] ^ input_a[7]);
  assign cgp_core_022 = ~(input_a[7] | input_a[2]);
  assign cgp_core_023 = ~(input_a[10] | input_a[5]);
  assign cgp_core_024 = input_a[2] ^ input_a[12];
  assign cgp_core_026 = input_a[11] & input_a[0];
  assign cgp_core_027 = ~input_a[3];
  assign cgp_core_030 = input_a[2] | input_a[4];
  assign cgp_core_031 = ~(input_a[5] | input_a[2]);
  assign cgp_core_032 = ~(input_a[6] & input_a[4]);
  assign cgp_core_033 = input_a[8] & input_a[8];
  assign cgp_core_034 = input_a[6] & input_a[0];
  assign cgp_core_036 = ~(input_a[8] | input_a[11]);
  assign cgp_core_038 = ~(input_a[6] & input_a[11]);
  assign cgp_core_039 = input_a[13] & input_a[0];
  assign cgp_core_041 = ~input_a[0];
  assign cgp_core_043 = ~(input_a[7] & input_a[3]);
  assign cgp_core_044 = ~(input_a[1] & input_a[0]);
  assign cgp_core_053 = ~input_a[10];
  assign cgp_core_054 = ~(input_a[1] & input_a[10]);
  assign cgp_core_056 = input_a[5] ^ input_a[4];
  assign cgp_core_057 = input_a[13] & input_a[10];
  assign cgp_core_058 = ~(input_a[6] | input_a[12]);
  assign cgp_core_060 = ~(input_a[8] | input_a[2]);
  assign cgp_core_061 = input_a[2] | input_a[7];
  assign cgp_core_062 = ~(input_a[9] & input_a[2]);
  assign cgp_core_063 = input_a[12] & input_a[8];
  assign cgp_core_066 = input_a[10] | input_a[8];
  assign cgp_core_067 = ~(input_a[4] & input_a[11]);
  assign cgp_core_069 = input_a[1] | input_a[0];
  assign cgp_core_070 = ~(input_a[6] ^ input_a[6]);
  assign cgp_core_071 = ~(input_a[11] | input_a[1]);
  assign cgp_core_076 = ~(input_a[12] | input_a[2]);
  assign cgp_core_077 = ~(input_a[4] ^ input_a[8]);
  assign cgp_core_078 = ~(input_a[12] | input_a[11]);
  assign cgp_core_080 = input_a[6] | input_a[7];
  assign cgp_core_081 = ~input_a[9];
  assign cgp_core_083 = ~(input_a[6] ^ input_a[4]);
  assign cgp_core_084 = input_a[9] ^ input_a[8];
  assign cgp_core_088 = ~(input_a[3] & input_a[1]);
  assign cgp_core_089 = ~(input_a[5] | input_a[3]);

  assign cgp_out[0] = input_a[9];
  assign cgp_out[1] = 1'b0;
  assign cgp_out[2] = 1'b0;
  assign cgp_out[3] = 1'b1;
endmodule