module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046_not;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_055_not;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_078;

  assign cgp_core_016 = input_f[1] ^ input_c[1];
  assign cgp_core_017 = input_c[0] & input_e[0];
  assign cgp_core_018 = ~(input_f[0] | input_e[1]);
  assign cgp_core_021 = input_f[0] & input_b[0];
  assign cgp_core_022 = input_a[0] | cgp_core_021;
  assign cgp_core_025 = ~(input_a[1] | input_a[1]);
  assign cgp_core_026 = ~(input_f[1] & input_f[1]);
  assign cgp_core_027 = ~input_g[1];
  assign cgp_core_029 = ~(input_a[0] & input_d[0]);
  assign cgp_core_030 = input_e[0] ^ cgp_core_029;
  assign cgp_core_031 = ~input_e[0];
  assign cgp_core_032 = ~input_b[0];
  assign cgp_core_033 = ~(input_g[0] | input_a[0]);
  assign cgp_core_036 = input_e[1] ^ cgp_core_033;
  assign cgp_core_037 = input_a[0] & input_b[0];
  assign cgp_core_039 = input_b[0] & input_e[0];
  assign cgp_core_040 = ~(input_g[1] & input_b[0]);
  assign cgp_core_041 = input_f[1] ^ input_c[1];
  assign cgp_core_042 = input_c[0] & input_e[1];
  assign cgp_core_043 = ~(cgp_core_041 & input_g[1]);
  assign cgp_core_044 = cgp_core_041 & input_a[0];
  assign cgp_core_046_not = ~cgp_core_039;
  assign cgp_core_047 = cgp_core_032 & cgp_core_039;
  assign cgp_core_048 = cgp_core_036 ^ cgp_core_043;
  assign cgp_core_049 = input_a[1] & cgp_core_043;
  assign cgp_core_055_not = ~input_e[0];
  assign cgp_core_060 = ~cgp_core_031;
  assign cgp_core_062 = ~(input_g[0] ^ input_g[0]);
  assign cgp_core_063 = input_d[1] & input_a[1];
  assign cgp_core_064 = ~(input_e[1] & input_f[0]);
  assign cgp_core_065 = input_d[1] & cgp_core_060;
  assign cgp_core_068 = input_c[0] & input_b[0];
  assign cgp_core_071 = input_b[0] ^ cgp_core_046_not;
  assign cgp_core_072 = input_f[1] & cgp_core_071;
  assign cgp_core_075 = input_g[0] | input_c[0];
  assign cgp_core_078 = ~input_e[1];

  assign cgp_out[0] = input_a[1];
endmodule