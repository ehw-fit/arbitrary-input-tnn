module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_015_not;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;

  assign cgp_core_015_not = ~input_c[0];
  assign cgp_core_016 = ~(input_d[1] & input_d[1]);
  assign cgp_core_017 = input_a[1] & input_a[1];
  assign cgp_core_018 = ~(input_c[2] & cgp_core_015_not);
  assign cgp_core_020 = input_b[2] ^ input_c[2];
  assign cgp_core_023 = input_d[0] & input_d[0];
  assign cgp_core_024 = ~input_d[1];
  assign cgp_core_025 = ~(input_b[1] ^ input_c[2]);
  assign cgp_core_026 = input_c[1] ^ input_d[0];
  assign cgp_core_029 = input_a[0] & input_b[2];
  assign cgp_core_030 = input_d[0] ^ input_c[0];
  assign cgp_core_031 = ~input_b[1];
  assign cgp_core_032 = ~(input_b[2] & input_a[1]);
  assign cgp_core_033 = input_c[2] ^ input_d[2];
  assign cgp_core_034 = input_a[1] ^ input_a[0];
  assign cgp_core_036 = ~(input_b[0] & input_d[2]);
  assign cgp_core_037 = ~(input_d[2] ^ input_a[1]);
  assign cgp_core_039 = input_b[2] & input_a[1];
  assign cgp_core_040 = input_b[2] ^ input_d[0];
  assign cgp_core_041 = ~input_b[1];
  assign cgp_core_042 = ~(input_c[2] & input_c[0]);
  assign cgp_core_044 = ~(input_b[2] ^ input_b[2]);
  assign cgp_core_046 = input_b[1] ^ cgp_core_030;
  assign cgp_core_047 = ~input_a[1];
  assign cgp_core_052 = input_b[1] | input_c[1];
  assign cgp_core_054 = ~(input_b[1] | input_d[0]);
  assign cgp_core_055 = input_d[1] | input_d[2];
  assign cgp_core_057 = ~(cgp_core_039 & input_d[2]);

  assign cgp_out[0] = input_b[2];
endmodule