module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = input_c[0] ^ input_d[0];
  assign cgp_core_017 = input_c[0] & input_d[0];
  assign cgp_core_018 = input_c[1] ^ input_d[1];
  assign cgp_core_019 = input_c[1] & input_d[1];
  assign cgp_core_020 = cgp_core_018 ^ cgp_core_017;
  assign cgp_core_021 = cgp_core_018 & cgp_core_017;
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_023 = input_e[0] ^ input_g[0];
  assign cgp_core_024 = input_e[0] & input_g[0];
  assign cgp_core_025 = input_e[1] ^ input_g[1];
  assign cgp_core_026 = input_e[1] & input_g[1];
  assign cgp_core_027 = cgp_core_025 ^ cgp_core_024;
  assign cgp_core_028 = cgp_core_025 & cgp_core_024;
  assign cgp_core_029 = cgp_core_026 | cgp_core_028;
  assign cgp_core_030 = cgp_core_016 ^ cgp_core_023;
  assign cgp_core_031 = cgp_core_016 & cgp_core_023;
  assign cgp_core_032 = cgp_core_020 ^ cgp_core_027;
  assign cgp_core_033 = cgp_core_020 & cgp_core_027;
  assign cgp_core_034 = cgp_core_032 ^ cgp_core_031;
  assign cgp_core_035 = cgp_core_032 & cgp_core_031;
  assign cgp_core_036 = cgp_core_033 | cgp_core_035;
  assign cgp_core_037 = cgp_core_022 ^ cgp_core_029;
  assign cgp_core_038 = cgp_core_022 & cgp_core_029;
  assign cgp_core_039 = cgp_core_037 ^ cgp_core_036;
  assign cgp_core_040 = cgp_core_037 & cgp_core_036;
  assign cgp_core_041 = cgp_core_038 | cgp_core_040;
  assign cgp_core_042 = input_b[0] ^ input_f[0];
  assign cgp_core_043 = input_b[0] & input_f[0];
  assign cgp_core_044 = input_b[1] ^ input_f[1];
  assign cgp_core_045 = input_b[1] & input_f[1];
  assign cgp_core_046 = cgp_core_044 ^ cgp_core_043;
  assign cgp_core_047 = cgp_core_044 & cgp_core_043;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = input_a[0] & cgp_core_042;
  assign cgp_core_051 = input_a[1] ^ cgp_core_046;
  assign cgp_core_052 = input_a[1] & cgp_core_046;
  assign cgp_core_053 = cgp_core_051 ^ cgp_core_050;
  assign cgp_core_054 = cgp_core_051 & cgp_core_050;
  assign cgp_core_055 = cgp_core_052 | cgp_core_054;
  assign cgp_core_056 = cgp_core_048 ^ cgp_core_055;
  assign cgp_core_057 = cgp_core_048 & cgp_core_055;
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = cgp_core_041 & cgp_core_058;
  assign cgp_core_060 = ~(cgp_core_041 ^ cgp_core_057);
  assign cgp_core_061 = ~cgp_core_056;
  assign cgp_core_062 = cgp_core_039 & cgp_core_061;
  assign cgp_core_063 = cgp_core_062 & cgp_core_060;
  assign cgp_core_064 = ~(cgp_core_039 ^ cgp_core_056);
  assign cgp_core_065 = cgp_core_064 & cgp_core_060;
  assign cgp_core_066 = ~cgp_core_053;
  assign cgp_core_067 = cgp_core_034 & cgp_core_066;
  assign cgp_core_068 = cgp_core_067 & cgp_core_065;
  assign cgp_core_069 = ~(cgp_core_034 ^ cgp_core_053);
  assign cgp_core_070 = cgp_core_069 & cgp_core_065;
  assign cgp_core_071 = input_f[0] ^ input_a[1];
  assign cgp_core_072 = ~(input_b[1] & input_e[0]);
  assign cgp_core_073 = input_e[0] ^ input_c[0];
  assign cgp_core_075 = cgp_core_030 & cgp_core_070;
  assign cgp_core_077 = cgp_core_059 | cgp_core_075;
  assign cgp_core_078 = cgp_core_063 | cgp_core_077;
  assign cgp_core_079 = cgp_core_068 | cgp_core_078;

  assign cgp_out[0] = cgp_core_079;
endmodule