module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_a[2] & input_a[2]);
  assign cgp_core_019 = ~input_b[1];
  assign cgp_core_024 = input_c[2] | input_d[2];
  assign cgp_core_026 = input_e[0] ^ input_b[0];
  assign cgp_core_027 = ~input_b[0];
  assign cgp_core_028 = ~input_c[1];
  assign cgp_core_030 = ~(input_c[1] | input_b[0]);
  assign cgp_core_034 = ~(input_e[1] & input_b[1]);
  assign cgp_core_036 = ~(input_c[0] & input_c[2]);
  assign cgp_core_038 = ~input_c[2];
  assign cgp_core_040 = input_e[0] & input_d[1];
  assign cgp_core_041 = input_e[2] ^ input_b[2];
  assign cgp_core_042 = ~input_c[2];
  assign cgp_core_044 = input_d[2] | input_e[1];
  assign cgp_core_046_not = ~input_b[1];
  assign cgp_core_049 = ~(input_c[2] | input_e[2]);
  assign cgp_core_050 = ~(input_a[1] | input_e[1]);
  assign cgp_core_051 = input_c[0] & input_d[1];
  assign cgp_core_058 = input_e[2] | input_b[0];
  assign cgp_core_059 = ~input_b[1];
  assign cgp_core_060 = input_a[2] & input_b[1];
  assign cgp_core_061 = ~(input_b[1] | input_b[1]);
  assign cgp_core_063 = ~(input_d[2] | input_d[2]);
  assign cgp_core_064 = ~(input_e[1] & input_c[2]);
  assign cgp_core_065 = ~(input_a[2] | input_a[2]);
  assign cgp_core_067 = ~(input_c[2] | input_d[0]);
  assign cgp_core_068 = ~input_e[1];
  assign cgp_core_070 = ~(input_d[2] & input_e[1]);
  assign cgp_core_072 = ~(input_b[2] & input_b[2]);
  assign cgp_core_076 = ~input_d[0];
  assign cgp_core_078 = ~(input_d[1] ^ input_c[0]);
  assign cgp_core_079 = input_c[1] ^ input_c[2];

  assign cgp_out[0] = cgp_core_049;
endmodule