module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_080;

  assign cgp_core_018 = ~(input_b[2] ^ input_b[1]);
  assign cgp_core_019 = ~(input_d[2] | input_e[1]);
  assign cgp_core_020 = ~(input_c[0] & input_c[1]);
  assign cgp_core_023 = ~(input_e[2] & input_c[1]);
  assign cgp_core_025 = ~input_a[0];
  assign cgp_core_027 = input_c[0] | input_c[2];
  assign cgp_core_033 = input_d[2] & input_d[2];
  assign cgp_core_034 = ~input_d[2];
  assign cgp_core_036 = ~(input_b[0] | input_c[0]);
  assign cgp_core_037 = input_a[2] ^ input_b[0];
  assign cgp_core_038 = ~(input_d[0] & input_a[1]);
  assign cgp_core_039 = ~input_e[1];
  assign cgp_core_040 = input_c[2] & input_d[0];
  assign cgp_core_041 = input_a[2] & input_a[1];
  assign cgp_core_044 = input_b[0] & input_c[0];
  assign cgp_core_046 = input_d[1] ^ input_c[0];
  assign cgp_core_047 = ~(input_e[2] & input_b[2]);
  assign cgp_core_049 = input_d[1] | input_c[1];
  assign cgp_core_050 = ~(input_b[0] ^ input_d[0]);
  assign cgp_core_051 = input_d[2] | input_b[1];
  assign cgp_core_052 = ~(input_a[1] & input_c[0]);
  assign cgp_core_053 = input_d[2] | input_c[2];
  assign cgp_core_054 = ~(input_b[0] & input_a[2]);
  assign cgp_core_056 = ~input_e[2];
  assign cgp_core_057 = ~cgp_core_053;
  assign cgp_core_058 = input_a[2] & cgp_core_057;
  assign cgp_core_060 = ~(input_a[2] ^ cgp_core_053);
  assign cgp_core_061 = cgp_core_060 & cgp_core_056;
  assign cgp_core_063 = ~input_c[0];
  assign cgp_core_064 = input_b[2] & cgp_core_061;
  assign cgp_core_067 = input_b[0] | input_d[0];
  assign cgp_core_068 = input_e[0] | input_d[0];
  assign cgp_core_069 = ~input_d[1];
  assign cgp_core_070 = ~(input_b[2] | input_b[1]);
  assign cgp_core_072 = ~input_b[0];
  assign cgp_core_074 = ~(input_c[0] | input_c[1]);
  assign cgp_core_075 = ~(input_b[2] ^ input_e[1]);
  assign cgp_core_076 = ~(input_d[1] & input_e[2]);
  assign cgp_core_080 = cgp_core_064 | cgp_core_058;

  assign cgp_out[0] = cgp_core_080;
endmodule