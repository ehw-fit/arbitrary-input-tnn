module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066_not;
  wire cgp_core_067;
  wire cgp_core_068_not;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076_not;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_019 = ~input_a[2];
  assign cgp_core_020 = input_b[2] & input_e[2];
  assign cgp_core_021 = ~(input_b[1] ^ input_e[2]);
  assign cgp_core_022 = ~(input_c[0] ^ input_c[1]);
  assign cgp_core_023 = input_b[2] ^ input_d[2];
  assign cgp_core_024_not = ~input_d[0];
  assign cgp_core_025 = input_a[0] & input_e[0];
  assign cgp_core_028 = input_b[2] | input_c[2];
  assign cgp_core_029 = ~(input_d[0] | input_b[1]);
  assign cgp_core_030 = ~(input_d[1] | input_d[2]);
  assign cgp_core_034 = ~(input_e[1] | input_a[2]);
  assign cgp_core_036 = input_d[2] & input_b[0];
  assign cgp_core_037 = input_d[0] & input_e[1];
  assign cgp_core_038 = ~(input_d[1] & input_c[2]);
  assign cgp_core_040 = ~(input_e[1] & input_a[0]);
  assign cgp_core_044 = input_a[0] ^ input_d[2];
  assign cgp_core_048 = ~(input_e[2] | input_e[2]);
  assign cgp_core_049 = ~(input_d[0] & input_a[2]);
  assign cgp_core_050 = ~(input_e[0] | input_d[2]);
  assign cgp_core_051 = input_d[1] & input_c[1];
  assign cgp_core_052 = input_e[2] | cgp_core_051;
  assign cgp_core_055 = input_d[2] | cgp_core_052;
  assign cgp_core_056 = input_e[2] | input_a[2];
  assign cgp_core_059 = ~cgp_core_028;
  assign cgp_core_060 = input_e[0] | input_d[0];
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_062 = cgp_core_061 & cgp_core_059;
  assign cgp_core_063 = ~input_e[1];
  assign cgp_core_064 = input_a[2] & cgp_core_063;
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066_not = ~input_c[2];
  assign cgp_core_067 = input_a[2] & cgp_core_062;
  assign cgp_core_068_not = ~input_a[0];
  assign cgp_core_069_not = ~input_e[1];
  assign cgp_core_070 = input_a[1] & cgp_core_067;
  assign cgp_core_071 = ~input_c[2];
  assign cgp_core_072 = ~(input_b[2] ^ input_a[2]);
  assign cgp_core_073 = input_b[2] | input_b[0];
  assign cgp_core_074 = ~(input_a[1] ^ input_d[1]);
  assign cgp_core_076_not = ~input_e[1];
  assign cgp_core_077 = input_b[2] & input_a[0];
  assign cgp_core_078 = cgp_core_070 | cgp_core_065;
  assign cgp_core_079 = input_e[1] | input_e[0];
  assign cgp_core_080 = input_b[0] ^ input_d[2];

  assign cgp_out[0] = cgp_core_078;
endmodule