module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_021_not;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_080;

  assign cgp_core_017 = ~(input_e[0] ^ input_e[0]);
  assign cgp_core_018 = input_e[1] ^ input_a[0];
  assign cgp_core_021_not = ~input_d[0];
  assign cgp_core_022 = ~input_c[0];
  assign cgp_core_023 = input_e[1] ^ input_d[0];
  assign cgp_core_024 = input_e[2] | input_a[2];
  assign cgp_core_025 = input_c[2] ^ input_e[2];
  assign cgp_core_029 = input_e[1] & input_b[1];
  assign cgp_core_030 = ~(input_b[0] | input_b[1]);
  assign cgp_core_033 = input_a[2] ^ input_a[2];
  assign cgp_core_036 = input_b[0] | input_d[2];
  assign cgp_core_038 = input_e[2] & input_d[1];
  assign cgp_core_039 = input_b[2] & input_e[0];
  assign cgp_core_041 = input_e[1] ^ input_c[1];
  assign cgp_core_045 = input_b[2] | input_e[1];
  assign cgp_core_048 = ~input_d[1];
  assign cgp_core_049 = ~input_c[1];
  assign cgp_core_053 = input_e[2] | input_d[2];
  assign cgp_core_054 = input_e[2] & input_d[2];
  assign cgp_core_055 = ~(input_a[2] & input_e[0]);
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_057 = ~cgp_core_053;
  assign cgp_core_058 = input_b[2] & cgp_core_057;
  assign cgp_core_061 = input_a[2] & cgp_core_056;
  assign cgp_core_062 = ~input_c[2];
  assign cgp_core_063 = input_b[1] & cgp_core_062;
  assign cgp_core_064 = cgp_core_063 & cgp_core_061;
  assign cgp_core_065 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_066 = input_e[2] & input_b[2];
  assign cgp_core_067 = ~input_c[0];
  assign cgp_core_068 = ~(input_e[1] & input_b[2]);
  assign cgp_core_069 = ~input_e[1];
  assign cgp_core_072 = input_e[1] ^ input_b[0];
  assign cgp_core_073 = input_d[1] ^ input_c[2];
  assign cgp_core_074 = ~input_a[1];
  assign cgp_core_075 = input_c[2] ^ input_c[0];
  assign cgp_core_080 = cgp_core_064 | cgp_core_058;

  assign cgp_out[0] = cgp_core_080;
endmodule