module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035_not;
  wire cgp_core_037_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051_not;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_059;
  wire cgp_core_063;
  wire cgp_core_066;

  assign cgp_core_015 = input_a[0] & input_c[0];
  assign cgp_core_016 = input_a[1] | input_c[1];
  assign cgp_core_017 = input_a[1] & input_c[1];
  assign cgp_core_019 = cgp_core_016 & cgp_core_015;
  assign cgp_core_020 = cgp_core_017 | cgp_core_019;
  assign cgp_core_022 = ~(input_c[1] | input_d[1]);
  assign cgp_core_023 = input_b[1] | input_d[1];
  assign cgp_core_024 = input_b[1] & input_d[1];
  assign cgp_core_025_not = ~input_e[1];
  assign cgp_core_026 = cgp_core_023 & input_d[0];
  assign cgp_core_027 = cgp_core_024 | cgp_core_026;
  assign cgp_core_028 = input_f[0] & input_b[1];
  assign cgp_core_029 = ~(input_b[0] | input_e[1]);
  assign cgp_core_030 = ~input_f[0];
  assign cgp_core_031 = input_e[1] & input_f[1];
  assign cgp_core_032 = ~(input_d[1] ^ input_b[1]);
  assign cgp_core_033 = input_c[1] ^ input_b[1];
  assign cgp_core_035_not = ~input_d[0];
  assign cgp_core_037_not = ~input_e[1];
  assign cgp_core_038 = input_f[1] | input_e[1];
  assign cgp_core_039 = ~(input_a[0] & input_a[0]);
  assign cgp_core_040 = ~(input_f[0] & input_c[1]);
  assign cgp_core_042 = cgp_core_027 | cgp_core_031;
  assign cgp_core_043 = input_e[0] | input_e[1];
  assign cgp_core_045 = input_a[0] ^ input_b[0];
  assign cgp_core_046 = ~(input_f[1] | input_b[0]);
  assign cgp_core_048 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_049 = ~cgp_core_042;
  assign cgp_core_050 = cgp_core_020 & cgp_core_049;
  assign cgp_core_051_not = ~input_f[0];
  assign cgp_core_052 = input_e[0] ^ input_d[1];
  assign cgp_core_053 = ~input_f[0];
  assign cgp_core_054_not = ~input_a[1];
  assign cgp_core_055 = input_a[0] & input_a[0];
  assign cgp_core_059 = input_e[0] ^ input_c[0];
  assign cgp_core_063 = ~input_d[0];
  assign cgp_core_066 = input_e[0] | input_e[0];

  assign cgp_out[0] = cgp_core_050;
endmodule