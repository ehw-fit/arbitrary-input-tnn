module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_079;

  assign cgp_core_018 = ~input_c[0];
  assign cgp_core_019 = ~(input_e[1] | input_e[1]);
  assign cgp_core_020 = ~input_f[1];
  assign cgp_core_021 = ~(input_c[0] | input_e[0]);
  assign cgp_core_022 = input_b[1] ^ input_e[0];
  assign cgp_core_023 = input_b[0] | input_f[1];
  assign cgp_core_025 = ~(input_c[0] ^ input_e[1]);
  assign cgp_core_028 = ~input_d[1];
  assign cgp_core_030 = ~(input_f[0] & input_c[1]);
  assign cgp_core_031 = ~(input_c[0] & input_d[0]);
  assign cgp_core_034 = input_a[1] & input_f[1];
  assign cgp_core_035 = ~(input_g[1] & input_a[1]);
  assign cgp_core_036 = ~input_f[1];
  assign cgp_core_037 = ~input_g[1];
  assign cgp_core_038 = ~input_b[1];
  assign cgp_core_040 = ~(input_b[0] ^ input_b[0]);
  assign cgp_core_041 = input_e[0] | input_e[1];
  assign cgp_core_042_not = ~input_e[1];
  assign cgp_core_043 = ~(input_f[0] | input_c[1]);
  assign cgp_core_045 = input_g[1] | input_b[1];
  assign cgp_core_046 = ~(input_g[0] ^ input_f[1]);
  assign cgp_core_047 = input_e[0] ^ input_g[1];
  assign cgp_core_048 = input_f[1] & input_c[1];
  assign cgp_core_049 = ~(input_f[1] ^ input_f[1]);
  assign cgp_core_050 = input_c[1] | input_d[0];
  assign cgp_core_051 = ~input_g[0];
  assign cgp_core_052 = ~(input_d[0] ^ input_e[0]);
  assign cgp_core_053 = input_f[1] | cgp_core_045;
  assign cgp_core_054 = input_f[1] & input_b[1];
  assign cgp_core_059 = ~(input_g[0] & input_b[0]);
  assign cgp_core_060 = ~(input_c[1] | cgp_core_054);
  assign cgp_core_061 = ~cgp_core_053;
  assign cgp_core_062 = input_d[1] & cgp_core_061;
  assign cgp_core_064 = input_c[0] | input_a[1];
  assign cgp_core_065 = input_e[1] & cgp_core_060;
  assign cgp_core_067 = ~input_e[0];
  assign cgp_core_068 = input_a[1] & cgp_core_065;
  assign cgp_core_069 = ~(input_d[0] | input_c[0]);
  assign cgp_core_070 = input_a[1] | input_c[0];
  assign cgp_core_071 = ~(input_b[0] & input_b[1]);
  assign cgp_core_072 = input_b[0] | input_f[1];
  assign cgp_core_073 = ~input_a[1];
  assign cgp_core_079 = cgp_core_068 | cgp_core_062;

  assign cgp_out[0] = cgp_core_079;
endmodule