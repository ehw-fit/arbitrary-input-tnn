module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_047_not;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059_not;
  wire cgp_core_061;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;

  assign cgp_core_014 = input_a[0] & input_d[0];
  assign cgp_core_016 = ~(input_b[0] & input_d[0]);
  assign cgp_core_017 = input_f[1] | input_f[0];
  assign cgp_core_018 = ~(input_d[0] | input_c[0]);
  assign cgp_core_019 = input_e[0] | input_a[0];
  assign cgp_core_021 = ~input_a[1];
  assign cgp_core_022 = ~(input_a[1] & input_e[1]);
  assign cgp_core_026 = ~input_a[1];
  assign cgp_core_027 = input_e[1] | input_f[1];
  assign cgp_core_028 = input_f[0] | input_b[1];
  assign cgp_core_031 = ~(input_e[0] ^ input_f[1]);
  assign cgp_core_033 = input_b[1] ^ input_a[1];
  assign cgp_core_034 = input_b[1] & input_a[0];
  assign cgp_core_035 = cgp_core_027 | input_d[1];
  assign cgp_core_036_not = ~input_e[0];
  assign cgp_core_037 = ~(input_a[1] | input_b[0]);
  assign cgp_core_038 = input_a[0] ^ input_a[0];
  assign cgp_core_039 = input_b[1] ^ input_d[1];
  assign cgp_core_040 = input_e[1] & input_f[1];
  assign cgp_core_044 = input_d[0] | cgp_core_035;
  assign cgp_core_045_not = ~input_f[1];
  assign cgp_core_047_not = ~input_d[1];
  assign cgp_core_048 = input_f[0] & input_b[0];
  assign cgp_core_049 = ~input_b[0];
  assign cgp_core_050 = ~(input_b[0] | input_f[0]);
  assign cgp_core_053 = input_c[0] & input_c[1];
  assign cgp_core_056 = ~input_b[0];
  assign cgp_core_057 = input_d[0] ^ input_f[1];
  assign cgp_core_059_not = ~input_a[0];
  assign cgp_core_061 = input_e[1] & input_b[0];
  assign cgp_core_065 = ~input_b[1];
  assign cgp_core_066 = ~input_f[1];
  assign cgp_core_068 = input_a[1] | cgp_core_044;
  assign cgp_core_069 = cgp_core_065 | cgp_core_068;
  assign cgp_core_070 = input_f[0] | input_c[1];
  assign cgp_core_072 = cgp_core_069 | input_c[1];

  assign cgp_out[0] = cgp_core_072;
endmodule