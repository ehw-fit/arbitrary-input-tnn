module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017_not;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051_not;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_056_not;
  wire cgp_core_057_not;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;

  assign cgp_core_016 = ~(input_a[0] ^ input_a[10]);
  assign cgp_core_017_not = ~input_a[5];
  assign cgp_core_019 = input_a[11] ^ input_a[8];
  assign cgp_core_022 = ~(input_a[10] & input_a[4]);
  assign cgp_core_023 = input_a[6] | input_a[11];
  assign cgp_core_024 = ~input_a[11];
  assign cgp_core_025 = ~(input_a[4] | input_a[12]);
  assign cgp_core_028 = input_a[1] ^ input_a[7];
  assign cgp_core_030 = ~(input_a[2] | input_a[8]);
  assign cgp_core_033 = input_a[2] & input_a[13];
  assign cgp_core_035 = ~(input_a[6] | input_a[2]);
  assign cgp_core_036 = ~input_a[4];
  assign cgp_core_037_not = ~input_a[1];
  assign cgp_core_038 = ~(input_a[11] | input_a[1]);
  assign cgp_core_040 = ~(input_a[3] ^ input_a[2]);
  assign cgp_core_041 = ~(input_a[9] ^ input_a[8]);
  assign cgp_core_042 = input_a[13] ^ input_a[11];
  assign cgp_core_044 = ~(input_a[4] ^ input_a[11]);
  assign cgp_core_045 = ~input_a[2];
  assign cgp_core_048 = ~(input_a[4] & input_a[0]);
  assign cgp_core_049 = input_a[8] & input_a[2];
  assign cgp_core_050 = input_a[7] & input_a[11];
  assign cgp_core_051_not = ~input_a[12];
  assign cgp_core_052 = input_a[4] ^ input_a[10];
  assign cgp_core_054 = ~(input_a[1] & input_a[8]);
  assign cgp_core_056_not = ~input_a[4];
  assign cgp_core_057_not = ~input_a[3];
  assign cgp_core_058 = ~(input_a[3] | input_a[6]);
  assign cgp_core_059 = ~input_a[1];
  assign cgp_core_060 = input_a[9] | input_a[1];
  assign cgp_core_061 = ~input_a[1];
  assign cgp_core_065 = input_a[13] | input_a[13];
  assign cgp_core_066 = ~(input_a[13] & input_a[9]);
  assign cgp_core_068 = ~input_a[1];
  assign cgp_core_069 = input_a[11] ^ input_a[3];
  assign cgp_core_076 = input_a[4] | input_a[1];
  assign cgp_core_077 = input_a[12] ^ input_a[12];
  assign cgp_core_078 = ~input_a[6];
  assign cgp_core_079 = input_a[6] ^ input_a[7];
  assign cgp_core_082 = ~input_a[9];
  assign cgp_core_083 = input_a[1] | input_a[9];
  assign cgp_core_084 = input_a[10] ^ input_a[9];
  assign cgp_core_086 = ~input_a[4];
  assign cgp_core_088 = ~(input_a[12] | input_a[0]);
  assign cgp_core_089 = input_a[3] & input_a[1];
  assign cgp_core_090 = ~(input_a[0] & input_a[10]);

  assign cgp_out[0] = 1'b1;
  assign cgp_out[1] = input_a[9];
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = input_a[3];
endmodule