module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030_not;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;

  assign cgp_core_014 = ~(input_a[0] & input_b[1]);
  assign cgp_core_015 = input_a[0] & input_c[0];
  assign cgp_core_016 = input_a[1] | input_c[1];
  assign cgp_core_020 = ~(input_c[0] ^ input_a[1]);
  assign cgp_core_021 = input_b[0] ^ input_d[0];
  assign cgp_core_022 = input_b[0] & input_a[1];
  assign cgp_core_023 = input_b[1] ^ input_e[1];
  assign cgp_core_024 = input_b[1] ^ input_c[1];
  assign cgp_core_025 = ~(cgp_core_023 & input_d[1]);
  assign cgp_core_026 = input_e[1] & input_b[0];
  assign cgp_core_027 = ~cgp_core_024;
  assign cgp_core_028 = input_e[0] ^ input_f[0];
  assign cgp_core_029 = input_e[0] & input_b[1];
  assign cgp_core_030_not = ~input_e[1];
  assign cgp_core_031 = input_e[1] & input_b[0];
  assign cgp_core_032 = ~input_f[0];
  assign cgp_core_033 = cgp_core_030_not | input_a[1];
  assign cgp_core_034 = cgp_core_031 | cgp_core_033;
  assign cgp_core_035 = cgp_core_021 ^ cgp_core_028;
  assign cgp_core_036 = cgp_core_021 & cgp_core_028;
  assign cgp_core_037 = cgp_core_025 ^ input_d[0];
  assign cgp_core_038 = cgp_core_025 | cgp_core_032;
  assign cgp_core_041 = cgp_core_038 | cgp_core_036;
  assign cgp_core_042 = ~(input_e[0] & cgp_core_034);
  assign cgp_core_044 = ~input_f[0];
  assign cgp_core_048 = ~input_f[0];
  assign cgp_core_051 = ~(input_a[1] | cgp_core_048);
  assign cgp_core_052 = ~(cgp_core_020 ^ input_c[1]);
  assign cgp_core_053 = cgp_core_052 & cgp_core_048;
  assign cgp_core_054 = ~(input_b[1] | cgp_core_037);
  assign cgp_core_056 = cgp_core_054 & cgp_core_053;
  assign cgp_core_059 = ~input_e[0];
  assign cgp_core_060 = input_b[0] ^ input_d[1];
  assign cgp_core_061 = input_d[0] & input_f[0];
  assign cgp_core_063 = ~input_f[0];
  assign cgp_core_064 = cgp_core_061 | cgp_core_056;
  assign cgp_core_065 = input_e[1] & input_f[1];
  assign cgp_core_066 = cgp_core_064 | input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule