module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;

  assign cgp_core_014 = input_a[0] ^ input_c[0];
  assign cgp_core_015 = input_a[0] & input_c[0];
  assign cgp_core_016 = input_a[1] ^ input_c[1];
  assign cgp_core_018 = cgp_core_016 ^ cgp_core_015;
  assign cgp_core_019 = cgp_core_016 & cgp_core_015;
  assign cgp_core_022 = input_e[0] & input_f[0];
  assign cgp_core_024 = input_c[0] & input_f[1];
  assign cgp_core_028 = ~input_d[0];
  assign cgp_core_031 = input_d[1] & cgp_core_022;
  assign cgp_core_032 = input_f[0] ^ input_d[0];
  assign cgp_core_033 = input_f[0] & input_d[0];
  assign cgp_core_034 = input_a[0] | cgp_core_033;
  assign cgp_core_035 = input_b[1] ^ cgp_core_034;
  assign cgp_core_036 = ~input_e[1];
  assign cgp_core_037 = cgp_core_014 ^ cgp_core_028;
  assign cgp_core_038 = cgp_core_014 & cgp_core_028;
  assign cgp_core_039 = cgp_core_018 ^ cgp_core_032;
  assign cgp_core_040 = cgp_core_018 & cgp_core_032;
  assign cgp_core_041 = input_b[0] ^ cgp_core_038;
  assign cgp_core_042 = input_b[0] & cgp_core_038;
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;
  assign cgp_core_048 = ~(input_a[1] | input_f[1]);
  assign cgp_core_049 = cgp_core_036 ^ cgp_core_048;
  assign cgp_core_050 = cgp_core_036 & cgp_core_048;
  assign cgp_core_051 = ~cgp_core_050;
  assign cgp_core_052 = cgp_core_049 & cgp_core_051;
  assign cgp_core_053 = ~input_e[1];
  assign cgp_core_054 = cgp_core_053 & cgp_core_051;
  assign cgp_core_055 = cgp_core_043 & cgp_core_054;
  assign cgp_core_056 = ~input_b[1];
  assign cgp_core_057 = cgp_core_056 & cgp_core_054;
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_059 = cgp_core_041 & cgp_core_058;
  assign cgp_core_060 = cgp_core_059 & cgp_core_057;
  assign cgp_core_061 = ~(cgp_core_041 ^ input_b[1]);
  assign cgp_core_062 = input_e[1] & cgp_core_057;
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_064 = cgp_core_037 & cgp_core_063;
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066 = ~(input_b[1] ^ input_b[0]);
  assign cgp_core_067 = cgp_core_066 & input_f[0];
  assign cgp_core_068 = cgp_core_060 | input_f[1];

  assign cgp_out[0] = 1'b1;
endmodule