module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_017 = ~(input_c[0] & input_b[2]);
  assign cgp_core_018 = input_b[0] ^ input_d[2];
  assign cgp_core_020 = input_d[1] & input_e[1];
  assign cgp_core_021 = ~(input_b[1] | input_e[2]);
  assign cgp_core_022 = ~(input_c[2] & input_a[0]);
  assign cgp_core_024 = ~(input_a[0] ^ input_c[1]);
  assign cgp_core_025 = ~(input_e[0] | input_b[0]);
  assign cgp_core_026_not = ~input_d[0];
  assign cgp_core_027 = input_c[2] | input_d[0];
  assign cgp_core_028 = ~(input_e[0] ^ input_a[0]);
  assign cgp_core_029_not = ~input_c[2];
  assign cgp_core_036 = ~input_a[1];
  assign cgp_core_037 = input_c[1] ^ input_d[1];
  assign cgp_core_038 = ~(input_c[0] ^ input_a[1]);
  assign cgp_core_041 = input_b[2] | input_b[2];
  assign cgp_core_044 = ~(input_a[0] & input_b[1]);
  assign cgp_core_046 = ~(input_a[2] & input_d[2]);
  assign cgp_core_047 = ~input_d[1];
  assign cgp_core_050 = ~input_b[1];
  assign cgp_core_051 = input_c[2] | input_e[2];
  assign cgp_core_054 = input_e[0] ^ input_b[0];
  assign cgp_core_057 = ~(input_d[0] ^ input_d[2]);
  assign cgp_core_061 = ~(input_b[1] | input_d[1]);
  assign cgp_core_063 = input_a[0] | input_e[1];
  assign cgp_core_064 = input_d[1] ^ input_a[0];
  assign cgp_core_065 = ~input_c[0];
  assign cgp_core_067 = input_a[1] ^ input_b[2];
  assign cgp_core_069 = ~(input_d[2] & input_e[1]);
  assign cgp_core_070 = input_d[1] | input_a[1];
  assign cgp_core_071 = ~(input_d[0] | input_c[2]);
  assign cgp_core_073 = ~(input_c[1] | input_a[1]);
  assign cgp_core_076 = ~input_c[2];
  assign cgp_core_077 = ~(input_a[1] | input_e[0]);
  assign cgp_core_078 = input_d[2] & input_d[1];

  assign cgp_out[0] = cgp_core_046;
endmodule