module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_056_not;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066_not;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072_not;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = input_c[1] | input_f[1];
  assign cgp_core_017 = input_b[1] ^ input_c[1];
  assign cgp_core_019 = input_c[0] | input_d[1];
  assign cgp_core_020 = input_e[1] & input_g[0];
  assign cgp_core_021 = ~input_b[0];
  assign cgp_core_024 = ~(input_c[0] ^ input_d[0]);
  assign cgp_core_025 = ~(input_f[0] ^ input_g[1]);
  assign cgp_core_026 = ~input_f[1];
  assign cgp_core_028 = input_e[0] ^ input_b[1];
  assign cgp_core_030 = ~(input_e[1] ^ input_f[1]);
  assign cgp_core_031 = input_a[1] & input_d[1];
  assign cgp_core_034 = input_b[1] | input_c[1];
  assign cgp_core_035 = input_b[1] & input_c[1];
  assign cgp_core_037 = cgp_core_034 & input_g[1];
  assign cgp_core_038 = cgp_core_035 | cgp_core_037;
  assign cgp_core_042 = ~input_d[0];
  assign cgp_core_044 = input_c[1] & input_f[0];
  assign cgp_core_046 = input_g[1] | input_d[1];
  assign cgp_core_047 = ~(input_c[1] | input_d[0]);
  assign cgp_core_048 = ~(input_c[0] & input_e[1]);
  assign cgp_core_049 = ~input_a[0];
  assign cgp_core_050_not = ~input_g[1];
  assign cgp_core_051 = ~input_a[1];
  assign cgp_core_053 = cgp_core_038 | input_f[1];
  assign cgp_core_056_not = ~input_g[0];
  assign cgp_core_058 = ~cgp_core_038;
  assign cgp_core_059 = cgp_core_031 & cgp_core_058;
  assign cgp_core_060 = ~(input_d[1] ^ cgp_core_038);
  assign cgp_core_061 = ~cgp_core_053;
  assign cgp_core_062 = input_e[1] & cgp_core_061;
  assign cgp_core_064 = ~(input_f[1] | input_g[0]);
  assign cgp_core_065 = input_a[0] & cgp_core_060;
  assign cgp_core_066_not = ~input_g[1];
  assign cgp_core_067 = input_e[1] & input_a[1];
  assign cgp_core_068 = cgp_core_067 & cgp_core_065;
  assign cgp_core_069 = input_c[1] | input_b[1];
  assign cgp_core_070 = ~(input_d[0] & input_a[0]);
  assign cgp_core_071 = ~(input_b[0] & input_g[0]);
  assign cgp_core_072_not = ~input_e[0];
  assign cgp_core_074 = ~(input_c[0] & input_g[0]);
  assign cgp_core_075 = ~(input_e[1] & input_d[0]);
  assign cgp_core_078 = cgp_core_062 | cgp_core_059;
  assign cgp_core_079 = cgp_core_068 | cgp_core_078;

  assign cgp_out[0] = cgp_core_079;
endmodule