module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014_not;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_057_not;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_014_not = ~input_b[0];
  assign cgp_core_015 = input_b[0] | input_a[0];
  assign cgp_core_016 = input_a[0] | input_c[1];
  assign cgp_core_017_not = ~input_c[1];
  assign cgp_core_018 = input_b[1] | input_d[0];
  assign cgp_core_020 = ~(input_f[1] | input_c[0]);
  assign cgp_core_021 = input_e[0] ^ input_f[0];
  assign cgp_core_022 = input_e[0] & input_f[0];
  assign cgp_core_026_not = ~input_a[0];
  assign cgp_core_027 = ~input_e[1];
  assign cgp_core_028 = input_d[0] ^ cgp_core_021;
  assign cgp_core_029 = input_d[0] & cgp_core_021;
  assign cgp_core_030 = input_f[1] | cgp_core_022;
  assign cgp_core_032 = cgp_core_030 | cgp_core_029;
  assign cgp_core_033 = input_e[0] | input_c[1];
  assign cgp_core_034 = ~input_f[1];
  assign cgp_core_035_not = ~input_e[1];
  assign cgp_core_037 = input_d[0] & input_f[0];
  assign cgp_core_038 = input_b[0] & cgp_core_028;
  assign cgp_core_039 = input_c[1] | cgp_core_032;
  assign cgp_core_040 = input_a[0] & input_c[0];
  assign cgp_core_041 = cgp_core_039 | cgp_core_038;
  assign cgp_core_042 = cgp_core_039 & cgp_core_038;
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;
  assign cgp_core_046 = input_d[1] | cgp_core_043;
  assign cgp_core_049 = input_e[1] | input_f[1];
  assign cgp_core_050 = ~input_a[0];
  assign cgp_core_053_not = ~input_e[0];
  assign cgp_core_054 = input_b[0] & input_e[1];
  assign cgp_core_057_not = ~input_c[1];
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_059 = cgp_core_041 & cgp_core_058;
  assign cgp_core_061 = ~(cgp_core_041 ^ input_b[1]);
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_065 = cgp_core_063 & cgp_core_061;
  assign cgp_core_068 = cgp_core_059 | cgp_core_046;
  assign cgp_core_069 = cgp_core_065 | cgp_core_068;
  assign cgp_core_070 = input_c[1] | input_a[1];
  assign cgp_core_071 = cgp_core_049 | cgp_core_070;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;

  assign cgp_out[0] = cgp_core_072;
endmodule