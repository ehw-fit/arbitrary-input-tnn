module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067_not;
  wire cgp_core_068_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078_not;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_098;

  assign cgp_core_020 = ~input_a[0];
  assign cgp_core_021 = input_a[0] & input_b[0];
  assign cgp_core_022 = input_a[1] ^ input_b[1];
  assign cgp_core_023 = ~input_a[1];
  assign cgp_core_024 = cgp_core_022 ^ cgp_core_021;
  assign cgp_core_025 = cgp_core_022 & cgp_core_021;
  assign cgp_core_026 = cgp_core_023 | cgp_core_025;
  assign cgp_core_027 = input_a[2] ^ input_b[2];
  assign cgp_core_028 = input_a[2] & input_b[2];
  assign cgp_core_029 = cgp_core_027 ^ cgp_core_026;
  assign cgp_core_030 = cgp_core_027 & cgp_core_026;
  assign cgp_core_032 = input_c[0] ^ input_d[0];
  assign cgp_core_033 = input_c[0] & input_d[0];
  assign cgp_core_034 = input_c[1] ^ input_d[1];
  assign cgp_core_035 = input_c[1] & input_d[1];
  assign cgp_core_036 = cgp_core_034 ^ cgp_core_033;
  assign cgp_core_037 = cgp_core_034 & cgp_core_033;
  assign cgp_core_038 = cgp_core_035 | cgp_core_037;
  assign cgp_core_039 = input_c[2] ^ input_d[2];
  assign cgp_core_040 = input_c[2] & input_d[2];
  assign cgp_core_041 = cgp_core_039 ^ cgp_core_038;
  assign cgp_core_042 = cgp_core_039 & cgp_core_038;
  assign cgp_core_043 = cgp_core_040 | input_f[1];
  assign cgp_core_044 = input_e[0] ^ input_f[0];
  assign cgp_core_047 = input_e[1] & input_f[1];
  assign cgp_core_051 = input_e[2] ^ input_f[2];
  assign cgp_core_052 = input_e[2] & input_d[1];
  assign cgp_core_056 = cgp_core_032 ^ cgp_core_044;
  assign cgp_core_057 = input_d[2] & cgp_core_044;
  assign cgp_core_062 = cgp_core_036 | input_f[1];
  assign cgp_core_063 = cgp_core_041 ^ cgp_core_051;
  assign cgp_core_064 = cgp_core_041 & cgp_core_051;
  assign cgp_core_065 = cgp_core_063 ^ cgp_core_062;
  assign cgp_core_067_not = ~cgp_core_064;
  assign cgp_core_068_not = ~cgp_core_043;
  assign cgp_core_070 = ~cgp_core_068_not;
  assign cgp_core_071 = cgp_core_068_not & cgp_core_067_not;
  assign cgp_core_072 = cgp_core_043 | cgp_core_071;
  assign cgp_core_073 = ~cgp_core_072;
  assign cgp_core_074 = ~cgp_core_072;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_078_not = ~cgp_core_070;
  assign cgp_core_079 = cgp_core_078_not & cgp_core_074;
  assign cgp_core_080 = ~cgp_core_065;
  assign cgp_core_085 = ~cgp_core_057;
  assign cgp_core_086 = cgp_core_024 & cgp_core_085;
  assign cgp_core_087 = cgp_core_086 & cgp_core_079;
  assign cgp_core_088 = ~(cgp_core_024 ^ cgp_core_057);
  assign cgp_core_089 = cgp_core_088 & cgp_core_079;
  assign cgp_core_093 = ~(cgp_core_020 ^ cgp_core_056);
  assign cgp_core_094 = cgp_core_093 & cgp_core_089;
  assign cgp_core_098 = cgp_core_087 | cgp_core_094;

  assign cgp_out[0] = 1'b0;
endmodule