module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018_not;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;

  assign cgp_core_017 = input_c[1] ^ input_c[0];
  assign cgp_core_018_not = ~input_c[1];
  assign cgp_core_019 = input_a[0] & input_b[2];
  assign cgp_core_020 = input_b[1] | input_c[1];
  assign cgp_core_022 = input_b[2] & input_d[1];
  assign cgp_core_023 = cgp_core_020 | cgp_core_022;
  assign cgp_core_029 = ~input_d[2];
  assign cgp_core_030 = ~input_c[2];
  assign cgp_core_031 = input_c[1] ^ input_e[1];
  assign cgp_core_032 = input_e[1] & input_e[1];
  assign cgp_core_033 = cgp_core_031 & cgp_core_030;
  assign cgp_core_034 = input_e[1] & cgp_core_030;
  assign cgp_core_035_not = ~input_c[1];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_041 = cgp_core_017 ^ cgp_core_029;
  assign cgp_core_042 = cgp_core_017 ^ input_d[1];
  assign cgp_core_044 = input_b[2] & cgp_core_033;
  assign cgp_core_046 = ~(input_c[2] | input_d[0]);
  assign cgp_core_047 = ~cgp_core_044;
  assign cgp_core_050 = ~input_a[2];
  assign cgp_core_051 = input_b[0] | cgp_core_047;
  assign cgp_core_052 = input_b[1] & input_b[2];
  assign cgp_core_054 = input_b[2] ^ input_e[0];
  assign cgp_core_055 = ~(input_d[0] | cgp_core_052);
  assign cgp_core_056 = ~(input_d[0] | cgp_core_052);
  assign cgp_core_057 = ~(cgp_core_054 ^ input_d[1]);
  assign cgp_core_058 = ~(cgp_core_057 ^ cgp_core_057);
  assign cgp_core_059 = input_a[0] | cgp_core_057;
  assign cgp_core_060 = ~input_e[1];
  assign cgp_core_063 = ~(input_a[0] ^ cgp_core_050);
  assign cgp_core_064 = input_b[0] & cgp_core_063;
  assign cgp_core_071 = ~input_b[0];
  assign cgp_core_073 = ~cgp_core_041;
  assign cgp_core_074 = input_a[0] & cgp_core_073;
  assign cgp_core_076 = ~input_a[0];

  assign cgp_out[0] = 1'b0;
endmodule