module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_059;

  assign cgp_core_014 = input_b[1] ^ input_d[1];
  assign cgp_core_018 = input_d[2] ^ input_c[0];
  assign cgp_core_019 = input_a[1] & input_a[1];
  assign cgp_core_022 = ~input_d[0];
  assign cgp_core_023 = input_c[1] ^ input_d[1];
  assign cgp_core_024 = ~(input_b[2] & input_c[2]);
  assign cgp_core_025 = cgp_core_022 & cgp_core_024;
  assign cgp_core_028 = ~(input_c[1] | input_d[2]);
  assign cgp_core_030 = input_b[2] ^ input_b[2];
  assign cgp_core_033_not = ~input_a[2];
  assign cgp_core_034 = input_c[2] ^ input_d[2];
  assign cgp_core_035 = input_a[2] ^ input_a[2];
  assign cgp_core_036 = input_c[1] & input_c[0];
  assign cgp_core_037 = ~cgp_core_034;
  assign cgp_core_038 = ~cgp_core_037;
  assign cgp_core_040 = input_a[1] & input_b[2];
  assign cgp_core_042 = ~cgp_core_023;
  assign cgp_core_044 = ~(cgp_core_023 ^ input_b[2]);
  assign cgp_core_045 = input_a[2] ^ input_d[0];
  assign cgp_core_047 = input_b[0] & input_a[1];
  assign cgp_core_048 = ~(input_b[0] & input_c[2]);
  assign cgp_core_049_not = ~input_c[0];
  assign cgp_core_050 = ~(input_c[1] & input_d[2]);
  assign cgp_core_052 = input_a[1] & input_b[2];
  assign cgp_core_053 = ~(input_b[1] ^ cgp_core_050);
  assign cgp_core_054 = ~(cgp_core_014 ^ input_c[2]);
  assign cgp_core_059 = input_b[1] | input_d[2];

  assign cgp_out[0] = 1'b1;
endmodule