module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_098;

  assign cgp_core_020 = input_d[2] ^ input_c[1];
  assign cgp_core_021 = input_a[0] & input_b[0];
  assign cgp_core_023 = input_a[0] ^ input_f[2];
  assign cgp_core_024_not = ~input_e[0];
  assign cgp_core_026 = input_b[1] | input_d[1];
  assign cgp_core_027 = input_c[2] ^ input_d[0];
  assign cgp_core_028 = ~(input_a[2] & input_e[1]);
  assign cgp_core_029 = input_d[2] & input_e[2];
  assign cgp_core_030 = cgp_core_027 & input_a[0];
  assign cgp_core_032 = input_f[1] ^ input_c[1];
  assign cgp_core_033 = input_b[0] & input_f[2];
  assign cgp_core_035 = ~(input_a[2] | input_a[0]);
  assign cgp_core_037 = ~input_d[0];
  assign cgp_core_040 = input_c[2] & input_b[0];
  assign cgp_core_041 = input_c[2] ^ input_a[0];
  assign cgp_core_043 = input_b[0] | input_b[1];
  assign cgp_core_044 = input_b[2] & input_e[1];
  assign cgp_core_045 = input_e[0] & input_f[0];
  assign cgp_core_046 = ~(input_e[1] | input_c[1]);
  assign cgp_core_047 = input_c[2] & input_f[1];
  assign cgp_core_048 = cgp_core_046 & input_a[2];
  assign cgp_core_049 = input_a[1] ^ input_c[0];
  assign cgp_core_050 = ~(input_b[2] ^ cgp_core_049);
  assign cgp_core_051 = input_e[2] ^ input_d[1];
  assign cgp_core_052 = input_a[1] & input_f[2];
  assign cgp_core_054 = input_c[1] & cgp_core_050;
  assign cgp_core_055 = ~cgp_core_052;
  assign cgp_core_057 = cgp_core_032 ^ cgp_core_044;
  assign cgp_core_060 = input_d[0] ^ input_b[0];
  assign cgp_core_061 = input_f[2] | cgp_core_057;
  assign cgp_core_063 = ~(cgp_core_041 | input_f[2]);
  assign cgp_core_066 = input_a[2] ^ input_e[1];
  assign cgp_core_069 = cgp_core_043 & cgp_core_055;
  assign cgp_core_070 = input_d[0] | input_a[2];
  assign cgp_core_071 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_073 = ~(cgp_core_069 | cgp_core_069);
  assign cgp_core_074 = ~input_a[0];
  assign cgp_core_075 = ~input_d[1];
  assign cgp_core_076 = ~input_d[2];
  assign cgp_core_077 = input_e[1] ^ input_e[2];
  assign cgp_core_079 = input_c[2] & input_d[2];
  assign cgp_core_081 = input_b[1] & input_a[2];
  assign cgp_core_082 = input_e[2] ^ input_d[0];
  assign cgp_core_083 = input_c[2] | input_d[1];
  assign cgp_core_084 = input_b[1] & input_e[0];
  assign cgp_core_085 = ~input_f[1];
  assign cgp_core_086 = cgp_core_024_not | cgp_core_085;
  assign cgp_core_087 = input_c[2] & input_a[0];
  assign cgp_core_088 = ~(cgp_core_024_not ^ input_c[1]);
  assign cgp_core_089 = ~input_c[2];
  assign cgp_core_090 = ~input_d[2];
  assign cgp_core_091 = input_b[2] & input_a[2];
  assign cgp_core_092 = cgp_core_091 & input_c[1];
  assign cgp_core_093 = input_f[0] | input_c[2];
  assign cgp_core_094 = ~(input_b[0] ^ input_c[0]);
  assign cgp_core_095 = input_e[1] | input_c[0];
  assign cgp_core_098 = ~(input_e[2] | input_c[2]);

  assign cgp_out[0] = 1'b0;
endmodule