module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047_not;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_073_not;
  wire cgp_core_074;
  wire cgp_core_075_not;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017_not = ~input_e[0];
  assign cgp_core_018 = ~(input_a[2] & input_c[1]);
  assign cgp_core_021 = ~(input_a[2] | input_b[0]);
  assign cgp_core_025 = ~input_c[0];
  assign cgp_core_027 = input_c[0] & input_c[2];
  assign cgp_core_028 = input_c[2] | input_e[2];
  assign cgp_core_029 = ~(input_c[2] & input_a[0]);
  assign cgp_core_030 = ~input_d[1];
  assign cgp_core_033 = ~(input_e[1] & input_b[2]);
  assign cgp_core_036 = ~(input_a[1] | input_e[1]);
  assign cgp_core_039 = input_a[0] ^ input_b[0];
  assign cgp_core_040 = ~(input_d[1] | input_e[1]);
  assign cgp_core_041 = cgp_core_028 | input_b[2];
  assign cgp_core_042 = input_c[2] & input_b[2];
  assign cgp_core_043_not = ~input_a[2];
  assign cgp_core_044 = ~(input_a[1] & input_b[2]);
  assign cgp_core_045 = input_e[2] ^ input_c[1];
  assign cgp_core_047_not = ~input_c[0];
  assign cgp_core_049_not = ~input_c[1];
  assign cgp_core_050 = input_c[2] | input_a[2];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_052_not = ~input_e[1];
  assign cgp_core_056 = ~cgp_core_051;
  assign cgp_core_057 = cgp_core_041 & cgp_core_056;
  assign cgp_core_059 = ~(input_e[2] ^ input_a[2]);
  assign cgp_core_061 = ~input_a[0];
  assign cgp_core_062 = ~input_c[2];
  assign cgp_core_065 = input_b[1] & cgp_core_059;
  assign cgp_core_066 = input_e[1] & input_e[0];
  assign cgp_core_067 = input_e[1] ^ input_b[2];
  assign cgp_core_068 = input_c[1] & cgp_core_065;
  assign cgp_core_069 = input_b[0] & input_e[1];
  assign cgp_core_071 = input_b[0] & input_c[0];
  assign cgp_core_073_not = ~input_b[2];
  assign cgp_core_074 = ~(input_b[2] & input_d[2]);
  assign cgp_core_075_not = ~input_e[2];
  assign cgp_core_079 = cgp_core_057 | cgp_core_042;
  assign cgp_core_080 = cgp_core_068 | cgp_core_079;

  assign cgp_out[0] = cgp_core_080;
endmodule