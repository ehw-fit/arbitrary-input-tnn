module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084_not;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088_not;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_094;
  wire cgp_core_098;

  assign cgp_core_020 = input_d[2] & input_f[2];
  assign cgp_core_021 = ~(input_c[1] & input_c[0]);
  assign cgp_core_022 = input_a[2] | input_a[0];
  assign cgp_core_023 = ~input_a[0];
  assign cgp_core_024 = ~input_f[2];
  assign cgp_core_026 = input_b[1] ^ input_e[1];
  assign cgp_core_030 = input_f[2] ^ input_e[2];
  assign cgp_core_032 = ~(input_f[0] ^ input_e[2]);
  assign cgp_core_033 = input_f[2] | input_a[0];
  assign cgp_core_035 = ~(input_c[1] | input_c[0]);
  assign cgp_core_037 = input_f[2] ^ input_e[2];
  assign cgp_core_039 = input_c[2] | input_d[2];
  assign cgp_core_040 = input_c[2] & input_d[2];
  assign cgp_core_044 = ~(input_a[2] | input_b[0]);
  assign cgp_core_047 = ~(input_a[0] ^ input_a[2]);
  assign cgp_core_048 = input_d[0] | input_f[2];
  assign cgp_core_050 = input_d[1] & input_f[0];
  assign cgp_core_051 = input_e[2] | input_f[2];
  assign cgp_core_052 = input_e[2] & input_f[2];
  assign cgp_core_053 = cgp_core_051 | cgp_core_050;
  assign cgp_core_054 = ~(input_e[0] | input_f[2]);
  assign cgp_core_056 = ~(input_a[2] | input_a[2]);
  assign cgp_core_057 = ~(input_f[2] ^ input_c[2]);
  assign cgp_core_058 = input_f[0] | input_a[0];
  assign cgp_core_059 = input_f[2] ^ input_c[0];
  assign cgp_core_060 = ~(input_e[0] | input_a[0]);
  assign cgp_core_062 = input_c[2] ^ input_a[1];
  assign cgp_core_063 = cgp_core_039 ^ cgp_core_053;
  assign cgp_core_064 = ~input_b[1];
  assign cgp_core_065 = ~cgp_core_063;
  assign cgp_core_067 = input_c[2] | cgp_core_063;
  assign cgp_core_068 = cgp_core_040 | cgp_core_052;
  assign cgp_core_070 = input_d[2] | cgp_core_067;
  assign cgp_core_074 = ~cgp_core_068;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = input_b[2] & cgp_core_075;
  assign cgp_core_079 = input_a[2] & cgp_core_074;
  assign cgp_core_080 = ~cgp_core_065;
  assign cgp_core_081 = input_b[2] & cgp_core_080;
  assign cgp_core_082 = cgp_core_081 & cgp_core_079;
  assign cgp_core_084_not = ~input_f[1];
  assign cgp_core_085 = input_f[1] & input_b[2];
  assign cgp_core_086 = input_c[0] ^ input_d[1];
  assign cgp_core_087 = ~input_e[1];
  assign cgp_core_088_not = ~input_f[1];
  assign cgp_core_090 = ~(input_e[2] ^ input_b[1]);
  assign cgp_core_092 = input_b[1] & input_e[1];
  assign cgp_core_094 = ~(input_e[0] | input_c[2]);
  assign cgp_core_098 = cgp_core_082 | cgp_core_076;

  assign cgp_out[0] = cgp_core_098;
endmodule