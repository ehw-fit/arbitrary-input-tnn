module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049_not;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_080;

  assign cgp_core_017 = ~input_c[2];
  assign cgp_core_018 = ~(input_a[0] ^ input_c[0]);
  assign cgp_core_020 = ~input_d[1];
  assign cgp_core_021 = ~(input_e[1] ^ input_d[2]);
  assign cgp_core_022 = input_e[0] | input_c[0];
  assign cgp_core_023 = input_b[1] | input_a[1];
  assign cgp_core_024 = input_a[2] | input_b[2];
  assign cgp_core_025 = input_e[2] & input_d[1];
  assign cgp_core_026_not = ~input_a[2];
  assign cgp_core_027 = cgp_core_024 & cgp_core_023;
  assign cgp_core_028 = input_d[2] | cgp_core_027;
  assign cgp_core_030 = input_c[2] ^ input_c[2];
  assign cgp_core_032 = input_a[1] & input_d[1];
  assign cgp_core_033 = ~(input_a[2] | input_e[1]);
  assign cgp_core_035 = ~(input_b[0] ^ input_e[1]);
  assign cgp_core_036 = input_a[1] ^ input_b[1];
  assign cgp_core_038 = ~(input_e[1] & input_d[1]);
  assign cgp_core_039 = input_b[1] | input_e[2];
  assign cgp_core_040 = input_a[2] | input_c[2];
  assign cgp_core_041 = input_e[2] ^ input_b[1];
  assign cgp_core_043 = input_a[0] ^ input_c[0];
  assign cgp_core_044 = input_d[0] & input_a[2];
  assign cgp_core_046 = ~input_d[1];
  assign cgp_core_047 = input_e[2] ^ input_b[2];
  assign cgp_core_048 = ~(input_a[2] & cgp_core_038);
  assign cgp_core_049_not = ~input_b[1];
  assign cgp_core_052 = ~(input_d[1] ^ input_b[1]);
  assign cgp_core_053 = ~input_e[2];
  assign cgp_core_055 = ~(input_a[2] | input_d[0]);
  assign cgp_core_056 = ~input_d[2];
  assign cgp_core_057 = ~input_c[2];
  assign cgp_core_058 = cgp_core_028 & cgp_core_057;
  assign cgp_core_059 = cgp_core_058 & cgp_core_056;
  assign cgp_core_060 = input_b[2] & cgp_core_053;
  assign cgp_core_062 = ~cgp_core_048;
  assign cgp_core_063 = input_b[2] & cgp_core_062;
  assign cgp_core_064 = cgp_core_063 & cgp_core_060;
  assign cgp_core_065 = ~input_a[0];
  assign cgp_core_066 = ~input_a[2];
  assign cgp_core_067 = ~(input_d[2] & input_e[2]);
  assign cgp_core_068 = ~(input_a[1] | input_d[0]);
  assign cgp_core_070 = ~(input_a[2] | input_d[0]);
  assign cgp_core_080 = cgp_core_064 | cgp_core_059;

  assign cgp_out[0] = cgp_core_080;
endmodule