module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_014 = ~(input_b[0] | input_b[1]);
  assign cgp_core_015 = input_b[1] & input_d[1];
  assign cgp_core_016 = input_c[0] ^ input_d[1];
  assign cgp_core_017 = ~(input_b[0] ^ input_d[1]);
  assign cgp_core_021 = ~(input_d[0] ^ input_a[1]);
  assign cgp_core_022 = ~(input_a[1] ^ input_d[1]);
  assign cgp_core_023 = ~input_e[0];
  assign cgp_core_024 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_025 = ~(input_c[0] | input_c[0]);
  assign cgp_core_026 = ~input_c[1];
  assign cgp_core_027 = input_d[0] ^ input_b[0];
  assign cgp_core_028 = input_e[1] & input_a[1];
  assign cgp_core_029_not = ~input_e[1];
  assign cgp_core_030 = ~(input_d[1] & input_a[0]);
  assign cgp_core_031 = ~(input_a[1] & input_b[1]);
  assign cgp_core_032 = input_e[1] ^ input_e[0];
  assign cgp_core_033 = input_c[1] | input_a[1];
  assign cgp_core_034 = input_a[1] & input_e[1];
  assign cgp_core_036 = ~cgp_core_034;
  assign cgp_core_037 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_039 = cgp_core_015 & cgp_core_036;
  assign cgp_core_040 = ~(input_e[1] | cgp_core_033);
  assign cgp_core_043 = ~input_c[0];
  assign cgp_core_044 = input_d[1] & cgp_core_040;
  assign cgp_core_045 = ~(input_b[1] ^ input_a[0]);
  assign cgp_core_047 = input_c[1] | input_b[1];
  assign cgp_core_048 = input_b[0] & input_a[0];
  assign cgp_core_049 = input_c[0] ^ input_e[1];
  assign cgp_core_051 = input_b[1] & cgp_core_040;
  assign cgp_core_053 = cgp_core_039 | cgp_core_051;
  assign cgp_core_054 = cgp_core_044 | cgp_core_053;

  assign cgp_out[0] = cgp_core_054;
endmodule