module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_083;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_100;
  wire cgp_core_101;
  wire cgp_core_104;
  wire cgp_core_105;

  assign cgp_core_020 = input_h[0] ^ input_i[0];
  assign cgp_core_023 = input_f[0] & input_i[1];
  assign cgp_core_025 = input_i[0] & input_i[0];
  assign cgp_core_026 = cgp_core_023 | input_b[1];
  assign cgp_core_027 = input_d[0] ^ cgp_core_020;
  assign cgp_core_028 = input_d[0] & input_f[0];
  assign cgp_core_030 = input_f[0] & input_f[1];
  assign cgp_core_032 = input_f[1] | cgp_core_028;
  assign cgp_core_033 = ~(input_c[1] ^ input_d[1]);
  assign cgp_core_034 = ~(input_h[1] & input_h[1]);
  assign cgp_core_035 = cgp_core_026 & cgp_core_033;
  assign cgp_core_037 = ~(input_h[0] ^ input_c[0]);
  assign cgp_core_038 = ~(input_b[1] & input_c[1]);
  assign cgp_core_041 = cgp_core_038 & input_a[1];
  assign cgp_core_042 = ~(input_f[1] & input_e[0]);
  assign cgp_core_043 = ~input_a[0];
  assign cgp_core_045 = input_a[1] ^ input_e[0];
  assign cgp_core_046 = ~input_i[0];
  assign cgp_core_047 = input_a[0] & input_a[0];
  assign cgp_core_048 = input_g[1] ^ input_f[0];
  assign cgp_core_050_not = ~cgp_core_042;
  assign cgp_core_051 = input_f[1] | input_d[1];
  assign cgp_core_052 = ~input_f[0];
  assign cgp_core_053 = input_g[0] & input_h[0];
  assign cgp_core_054 = input_f[1] ^ input_i[0];
  assign cgp_core_056 = input_c[0] & input_i[1];
  assign cgp_core_057 = cgp_core_054 & input_c[0];
  assign cgp_core_058 = ~(input_d[1] & input_e[0]);
  assign cgp_core_059 = ~input_e[0];
  assign cgp_core_061 = input_e[1] ^ input_e[1];
  assign cgp_core_062 = ~(input_h[1] & input_i[0]);
  assign cgp_core_063 = input_c[0] ^ input_f[0];
  assign cgp_core_064 = input_e[1] & input_c[1];
  assign cgp_core_065 = cgp_core_062 & input_f[0];
  assign cgp_core_066 = cgp_core_058 ^ cgp_core_065;
  assign cgp_core_070 = cgp_core_047 | input_c[0];
  assign cgp_core_071 = cgp_core_047 & cgp_core_063;
  assign cgp_core_075 = ~(cgp_core_050_not & cgp_core_066);
  assign cgp_core_076 = cgp_core_050_not & input_f[0];
  assign cgp_core_077 = input_h[0] ^ input_e[1];
  assign cgp_core_079 = cgp_core_076 ^ input_d[1];
  assign cgp_core_080 = cgp_core_051 & input_c[0];
  assign cgp_core_083 = ~(cgp_core_080 & input_d[0]);
  assign cgp_core_086 = ~input_h[0];
  assign cgp_core_088 = ~(input_f[0] & input_g[0]);
  assign cgp_core_091 = input_c[0] & input_g[0];
  assign cgp_core_092 = ~input_i[0];
  assign cgp_core_093 = ~(input_h[0] ^ cgp_core_092);
  assign cgp_core_094 = cgp_core_093 | cgp_core_091;
  assign cgp_core_096 = input_h[0] & input_h[1];
  assign cgp_core_097 = ~input_h[0];
  assign cgp_core_100 = ~(input_f[1] ^ input_h[1]);
  assign cgp_core_101 = input_e[1] & input_b[1];
  assign cgp_core_104 = input_a[1] & cgp_core_101;
  assign cgp_core_105 = input_c[0] & input_g[0];

  assign cgp_out[0] = 1'b0;
endmodule