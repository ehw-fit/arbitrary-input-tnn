module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030_not;
  wire cgp_core_031;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;

  assign cgp_core_011 = ~input_b[0];
  assign cgp_core_012 = input_b[1] ^ input_c[1];
  assign cgp_core_014 = input_b[1] | input_b[1];
  assign cgp_core_015 = input_c[0] | input_b[0];
  assign cgp_core_016_not = ~input_c[1];
  assign cgp_core_017 = input_a[1] | input_a[1];
  assign cgp_core_020 = ~input_a[2];
  assign cgp_core_021 = input_b[1] | input_c[1];
  assign cgp_core_022 = input_c[2] | input_a[2];
  assign cgp_core_023 = input_a[1] ^ input_c[0];
  assign cgp_core_024 = ~cgp_core_022;
  assign cgp_core_025 = ~input_c[0];
  assign cgp_core_027 = input_b[2] & cgp_core_024;
  assign cgp_core_028 = ~(input_a[0] ^ input_c[2]);
  assign cgp_core_029 = input_b[2] ^ input_a[0];
  assign cgp_core_030_not = ~input_b[0];
  assign cgp_core_031 = input_c[2] ^ input_a[1];
  assign cgp_core_032_not = ~input_c[1];
  assign cgp_core_033 = ~(input_b[1] ^ input_b[2]);
  assign cgp_core_034_not = ~input_b[0];
  assign cgp_core_035 = input_c[0] & input_b[2];
  assign cgp_core_037 = ~(input_a[1] ^ input_c[0]);
  assign cgp_core_038_not = ~input_c[1];
  assign cgp_core_040 = input_b[0] | input_b[1];
  assign cgp_core_041 = input_b[0] ^ input_b[0];
  assign cgp_core_042 = input_b[2] | input_a[2];

  assign cgp_out[0] = cgp_core_027;
endmodule