module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_016_not = ~input_d[1];
  assign cgp_core_017 = input_d[1] & input_d[1];
  assign cgp_core_019 = ~(input_a[2] ^ input_a[1]);
  assign cgp_core_020 = input_b[1] | input_a[1];
  assign cgp_core_021 = input_a[2] | input_b[2];
  assign cgp_core_023 = cgp_core_021 | input_a[1];
  assign cgp_core_024 = cgp_core_021 & cgp_core_020;
  assign cgp_core_028 = input_d[1] | input_b[2];
  assign cgp_core_029 = input_c[1] & input_d[1];
  assign cgp_core_031 = input_c[2] & input_d[2];
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_033 = input_c[2] | input_d[2];
  assign cgp_core_034 = input_c[0] & input_b[1];
  assign cgp_core_035 = cgp_core_033 | cgp_core_032;
  assign cgp_core_036 = cgp_core_033 & cgp_core_032;
  assign cgp_core_038 = ~cgp_core_036;
  assign cgp_core_039 = cgp_core_024 & cgp_core_038;
  assign cgp_core_041 = ~cgp_core_035;
  assign cgp_core_042 = cgp_core_023 & cgp_core_041;
  assign cgp_core_044 = ~(input_b[1] ^ input_b[0]);
  assign cgp_core_045 = input_d[2] ^ input_d[1];
  assign cgp_core_048 = input_a[2] ^ input_c[1];
  assign cgp_core_049 = ~(input_b[2] & input_b[2]);
  assign cgp_core_050 = ~(input_b[2] ^ input_b[0]);
  assign cgp_core_052 = ~input_c[0];
  assign cgp_core_053 = input_d[0] ^ input_b[1];
  assign cgp_core_055 = input_a[2] & input_b[2];
  assign cgp_core_057 = cgp_core_039 | cgp_core_055;
  assign cgp_core_058 = cgp_core_042 | cgp_core_057;
  assign cgp_core_059 = input_c[2] | input_b[0];

  assign cgp_out[0] = cgp_core_058;
endmodule