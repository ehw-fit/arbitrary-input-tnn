module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015_not;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046_not;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056_not;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059_not;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_069;

  assign cgp_core_014 = input_a[0] & input_d[0];
  assign cgp_core_015_not = ~input_d[1];
  assign cgp_core_016 = input_a[1] & input_b[1];
  assign cgp_core_017 = input_d[0] & input_c[1];
  assign cgp_core_018 = ~(input_b[1] & cgp_core_015_not);
  assign cgp_core_022 = ~(input_d[0] ^ input_d[0]);
  assign cgp_core_023 = input_f[1] | input_f[1];
  assign cgp_core_024 = ~(input_d[1] & input_e[0]);
  assign cgp_core_025 = ~(cgp_core_023 ^ input_f[0]);
  assign cgp_core_026 = input_e[0] & input_c[0];
  assign cgp_core_028 = ~(input_d[1] ^ input_d[0]);
  assign cgp_core_029_not = ~input_a[1];
  assign cgp_core_033 = input_e[1] & cgp_core_029_not;
  assign cgp_core_034 = ~input_d[1];
  assign cgp_core_039 = input_f[0] ^ input_d[1];
  assign cgp_core_041 = ~input_c[0];
  assign cgp_core_042 = input_d[0] & input_b[0];
  assign cgp_core_043 = ~input_b[1];
  assign cgp_core_044 = input_e[0] ^ input_e[0];
  assign cgp_core_045 = input_d[0] ^ input_e[0];
  assign cgp_core_046_not = ~input_f[0];
  assign cgp_core_047 = ~input_c[0];
  assign cgp_core_048 = input_b[0] | input_c[0];
  assign cgp_core_051 = ~input_e[1];
  assign cgp_core_052 = ~(input_b[0] & cgp_core_051);
  assign cgp_core_055 = ~input_a[0];
  assign cgp_core_056_not = ~input_b[0];
  assign cgp_core_057 = ~(input_e[0] | input_b[0]);
  assign cgp_core_058 = ~(input_a[1] & input_b[1]);
  assign cgp_core_059_not = ~input_e[1];
  assign cgp_core_060 = cgp_core_059_not & cgp_core_057;
  assign cgp_core_061 = input_f[1] | input_d[0];
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_069 = ~(input_b[1] | input_c[1]);

  assign cgp_out[0] = 1'b1;
endmodule