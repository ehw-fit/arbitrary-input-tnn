module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_013;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_026_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;

  assign cgp_core_013 = input_b[1] ^ input_b[1];
  assign cgp_core_015 = input_a[0] ^ input_d[1];
  assign cgp_core_017 = ~(input_e[1] | input_a[1]);
  assign cgp_core_019 = input_b[0] ^ input_a[0];
  assign cgp_core_020 = ~(input_b[0] | input_d[0]);
  assign cgp_core_021 = input_b[0] & input_a[1];
  assign cgp_core_026_not = ~input_b[0];
  assign cgp_core_028 = input_b[0] & input_a[0];
  assign cgp_core_029 = input_d[1] & input_d[0];
  assign cgp_core_034 = input_d[1] ^ input_b[1];
  assign cgp_core_036 = ~input_e[1];
  assign cgp_core_037_not = ~input_b[1];
  assign cgp_core_038 = input_e[0] & input_c[0];
  assign cgp_core_039 = input_d[0] | input_d[1];
  assign cgp_core_040 = ~input_a[1];
  assign cgp_core_041 = input_d[1] & input_e[1];
  assign cgp_core_042 = ~(input_b[0] | input_b[1]);
  assign cgp_core_043 = ~input_e[1];
  assign cgp_core_045 = input_d[1] ^ input_c[1];
  assign cgp_core_046 = ~(input_e[1] & input_a[0]);
  assign cgp_core_047 = input_e[0] ^ input_d[1];
  assign cgp_core_049 = ~input_a[1];
  assign cgp_core_050 = input_e[1] | input_d[1];
  assign cgp_core_051 = ~(input_d[1] ^ input_a[0]);
  assign cgp_core_052 = ~input_b[1];
  assign cgp_core_053 = input_e[1] ^ input_c[1];
  assign cgp_core_054 = ~input_c[0];

  assign cgp_out[0] = cgp_core_017;
endmodule