module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043_not;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;

  assign cgp_core_016 = ~(input_g[0] & input_c[0]);
  assign cgp_core_022 = ~(input_d[0] ^ input_e[1]);
  assign cgp_core_023 = ~input_a[0];
  assign cgp_core_024 = input_b[1] ^ input_a[0];
  assign cgp_core_025 = ~input_d[1];
  assign cgp_core_027 = cgp_core_025 & input_c[0];
  assign cgp_core_029 = ~input_d[0];
  assign cgp_core_030 = input_f[0] & input_c[1];
  assign cgp_core_031 = ~(input_d[0] | input_b[0]);
  assign cgp_core_032 = input_e[0] ^ input_c[1];
  assign cgp_core_033 = input_d[1] | input_d[1];
  assign cgp_core_034 = input_e[0] | input_f[1];
  assign cgp_core_035 = ~input_a[1];
  assign cgp_core_037 = cgp_core_034 & cgp_core_033;
  assign cgp_core_038 = input_e[1] & input_d[0];
  assign cgp_core_039 = input_f[1] ^ input_e[0];
  assign cgp_core_040 = input_g[1] & input_g[0];
  assign cgp_core_041 = ~(input_a[1] & input_g[1]);
  assign cgp_core_043_not = ~input_c[0];
  assign cgp_core_046 = ~input_c[0];
  assign cgp_core_049 = input_b[0] & input_e[1];
  assign cgp_core_053 = cgp_core_038 & input_g[0];
  assign cgp_core_054 = ~(input_f[0] ^ input_c[0]);
  assign cgp_core_055 = input_d[0] ^ input_f[0];
  assign cgp_core_057 = ~input_g[0];
  assign cgp_core_059 = input_c[0] & input_g[1];
  assign cgp_core_060 = input_b[1] & input_d[1];
  assign cgp_core_061 = input_e[1] & input_e[0];
  assign cgp_core_065 = input_c[1] & input_f[1];
  assign cgp_core_066 = input_e[1] & input_d[1];
  assign cgp_core_068 = input_a[1] & input_e[1];
  assign cgp_core_069 = input_f[1] & input_a[1];
  assign cgp_core_070 = cgp_core_069 & input_d[0];
  assign cgp_core_071 = ~(input_b[1] & cgp_core_046);
  assign cgp_core_073 = ~(input_f[1] & input_a[0]);
  assign cgp_core_074_not = ~input_g[1];
  assign cgp_core_075 = ~(cgp_core_074_not | input_c[0]);
  assign cgp_core_076 = cgp_core_073 | input_b[1];
  assign cgp_core_077 = input_a[1] & input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule