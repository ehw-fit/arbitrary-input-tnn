module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;

  assign cgp_core_017_not = ~input_e[0];
  assign cgp_core_018 = input_e[0] & input_e[0];
  assign cgp_core_020 = input_b[2] | input_b[2];
  assign cgp_core_023 = cgp_core_020 | input_a[1];
  assign cgp_core_026 = input_d[1] ^ input_a[0];
  assign cgp_core_028_not = ~input_e[2];
  assign cgp_core_029 = input_c[0] ^ input_e[1];
  assign cgp_core_030 = input_b[2] & cgp_core_017_not;
  assign cgp_core_032 = input_b[1] & input_d[1];
  assign cgp_core_033 = ~input_b[1];
  assign cgp_core_034 = input_b[1] & cgp_core_030;
  assign cgp_core_035 = cgp_core_032 | input_e[1];
  assign cgp_core_037 = ~(input_b[2] ^ cgp_core_026);
  assign cgp_core_039 = ~input_b[2];
  assign cgp_core_043 = input_a[0] ^ input_d[0];
  assign cgp_core_044 = input_d[2] & input_d[0];
  assign cgp_core_045 = ~(input_a[1] ^ input_c[2]);
  assign cgp_core_046 = input_c[2] & input_e[1];
  assign cgp_core_047 = input_a[2] ^ cgp_core_044;
  assign cgp_core_048 = input_c[1] | cgp_core_044;
  assign cgp_core_049 = cgp_core_046 | cgp_core_048;
  assign cgp_core_050 = input_a[2] ^ input_e[0];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_052 = cgp_core_050 ^ cgp_core_049;
  assign cgp_core_053 = cgp_core_050 & cgp_core_049;
  assign cgp_core_054 = input_e[1] | input_e[2];
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_057 = ~(input_c[2] & input_c[2]);
  assign cgp_core_069 = ~(input_a[0] ^ cgp_core_047);
  assign cgp_core_070 = cgp_core_069 & input_e[2];
  assign cgp_core_071 = ~input_a[2];
  assign cgp_core_073 = input_e[2] | input_a[0];
  assign cgp_core_074 = ~(input_e[2] | cgp_core_043);
  assign cgp_core_075 = ~cgp_core_074;

  assign cgp_out[0] = 1'b1;
endmodule