module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_068;

  assign cgp_core_014 = input_a[0] ^ input_c[0];
  assign cgp_core_015 = input_a[0] & input_c[0];
  assign cgp_core_016 = input_b[0] ^ input_c[1];
  assign cgp_core_017 = input_b[1] & input_c[0];
  assign cgp_core_018 = cgp_core_016 ^ input_f[1];
  assign cgp_core_019 = ~cgp_core_016;
  assign cgp_core_020 = cgp_core_017 | cgp_core_019;
  assign cgp_core_021 = input_e[0] ^ input_f[0];
  assign cgp_core_023 = input_e[1] | input_f[1];
  assign cgp_core_024 = ~input_e[1];
  assign cgp_core_026 = cgp_core_023 & input_f[0];
  assign cgp_core_028 = ~input_b[1];
  assign cgp_core_029 = ~input_d[0];
  assign cgp_core_037 = cgp_core_014 ^ cgp_core_028;
  assign cgp_core_038 = cgp_core_014 & cgp_core_028;
  assign cgp_core_041_not = ~input_b[0];
  assign cgp_core_042 = input_d[1] & input_e[1];
  assign cgp_core_043 = cgp_core_018 | cgp_core_042;
  assign cgp_core_044 = cgp_core_020 ^ input_e[0];
  assign cgp_core_045 = ~input_d[1];
  assign cgp_core_046 = cgp_core_044 ^ cgp_core_043;
  assign cgp_core_047 = cgp_core_044 | cgp_core_043;
  assign cgp_core_051 = ~input_a[1];
  assign cgp_core_054 = input_d[0] & cgp_core_051;
  assign cgp_core_055 = cgp_core_046 & cgp_core_054;
  assign cgp_core_056 = ~cgp_core_046;
  assign cgp_core_057 = cgp_core_056 & cgp_core_054;
  assign cgp_core_060 = ~cgp_core_041_not;
  assign cgp_core_061 = ~(cgp_core_041_not ^ input_b[1]);
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_064 = input_d[0] & cgp_core_063;
  assign cgp_core_068 = cgp_core_060 | cgp_core_055;

  assign cgp_out[0] = 1'b1;
endmodule