module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_027_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058_not;

  assign cgp_core_014 = ~input_c[1];
  assign cgp_core_017 = input_d[2] | input_b[1];
  assign cgp_core_020 = input_a[2] | input_a[1];
  assign cgp_core_022 = input_c[2] & input_a[2];
  assign cgp_core_023 = ~(input_a[0] ^ input_c[1]);
  assign cgp_core_024 = input_a[1] & input_c[0];
  assign cgp_core_025_not = ~input_c[2];
  assign cgp_core_027_not = ~input_a[1];
  assign cgp_core_028 = input_d[2] & input_a[1];
  assign cgp_core_029 = ~(input_a[1] | input_c[2]);
  assign cgp_core_030 = ~(input_d[1] | input_d[0]);
  assign cgp_core_031 = input_b[0] | input_a[2];
  assign cgp_core_034 = ~(input_c[2] | input_d[2]);
  assign cgp_core_036 = ~(input_d[0] & input_a[2]);
  assign cgp_core_038 = ~(input_c[0] ^ input_d[0]);
  assign cgp_core_039 = input_a[2] & input_b[1];
  assign cgp_core_040_not = ~input_b[2];
  assign cgp_core_041 = ~input_b[2];
  assign cgp_core_042 = ~(input_d[1] ^ input_a[2]);
  assign cgp_core_045 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_046 = ~input_b[2];
  assign cgp_core_047_not = ~input_a[1];
  assign cgp_core_049 = ~input_b[0];
  assign cgp_core_050 = input_c[0] ^ input_d[2];
  assign cgp_core_051 = ~(input_d[2] | input_c[2]);
  assign cgp_core_052 = ~cgp_core_014;
  assign cgp_core_053 = ~(input_d[1] ^ input_b[2]);
  assign cgp_core_054 = input_b[1] ^ input_c[0];
  assign cgp_core_055 = ~input_d[0];
  assign cgp_core_056 = ~input_d[1];
  assign cgp_core_057 = input_d[0] ^ input_a[0];
  assign cgp_core_058_not = ~input_b[2];

  assign cgp_out[0] = input_b[2];
endmodule