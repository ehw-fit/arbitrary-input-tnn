module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_011_not;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;

  assign cgp_core_011_not = ~input_a[2];
  assign cgp_core_012 = input_b[2] | input_c[1];
  assign cgp_core_013 = input_b[2] ^ input_a[2];
  assign cgp_core_014 = ~input_b[1];
  assign cgp_core_015 = ~(input_c[1] & input_a[0]);
  assign cgp_core_017 = input_b[2] & input_b[0];
  assign cgp_core_021 = input_c[0] | input_b[1];
  assign cgp_core_025 = input_b[0] ^ input_a[2];
  assign cgp_core_026 = ~input_b[2];
  assign cgp_core_027 = ~(input_c[0] & input_a[0]);
  assign cgp_core_029 = ~(input_c[0] ^ input_c[1]);
  assign cgp_core_030 = input_a[2] | input_b[1];
  assign cgp_core_031 = ~(input_b[1] & input_a[2]);
  assign cgp_core_033 = ~input_a[2];
  assign cgp_core_035 = input_c[2] & input_c[2];
  assign cgp_core_038 = input_a[0] ^ input_c[0];
  assign cgp_core_040 = ~(input_a[0] ^ input_c[0]);
  assign cgp_core_042 = ~(input_a[2] & input_a[2]);

  assign cgp_out[0] = 1'b1;
endmodule