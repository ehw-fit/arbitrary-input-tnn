module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030_not;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_056_not;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_070_not;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080_not;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_097;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_101;
  wire cgp_core_103;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_108;

  assign cgp_core_021 = ~(input_e[0] | input_c[1]);
  assign cgp_core_022 = ~(input_g[1] | input_d[0]);
  assign cgp_core_027 = input_i[0] ^ input_h[0];
  assign cgp_core_028 = input_c[0] | input_f[1];
  assign cgp_core_030_not = ~input_d[1];
  assign cgp_core_032 = ~(input_g[0] | input_i[0]);
  assign cgp_core_034 = input_f[0] ^ input_e[1];
  assign cgp_core_036 = ~input_c[0];
  assign cgp_core_039 = ~(input_g[0] ^ input_d[0]);
  assign cgp_core_042 = input_e[1] | input_d[1];
  assign cgp_core_043 = ~input_e[0];
  assign cgp_core_044 = input_c[1] & input_b[0];
  assign cgp_core_045 = input_a[1] | input_a[0];
  assign cgp_core_048 = input_c[1] ^ input_c[0];
  assign cgp_core_049 = input_f[0] & input_g[1];
  assign cgp_core_050 = ~input_i[1];
  assign cgp_core_051 = input_g[1] | input_e[0];
  assign cgp_core_052 = ~input_e[0];
  assign cgp_core_054 = input_h[1] | input_i[0];
  assign cgp_core_056_not = ~input_a[1];
  assign cgp_core_057 = input_e[1] & input_f[1];
  assign cgp_core_058 = ~input_g[1];
  assign cgp_core_059 = input_g[0] | input_e[0];
  assign cgp_core_061 = input_e[1] | input_g[1];
  assign cgp_core_062 = input_e[1] & input_g[1];
  assign cgp_core_064 = ~(input_c[0] | input_a[1]);
  assign cgp_core_066 = input_f[1] | cgp_core_062;
  assign cgp_core_067 = ~(input_i[1] | input_d[1]);
  assign cgp_core_068 = ~(input_g[1] | input_h[1]);
  assign cgp_core_069_not = ~input_g[0];
  assign cgp_core_070_not = ~input_d[1];
  assign cgp_core_071 = cgp_core_045 & cgp_core_061;
  assign cgp_core_072 = input_f[0] ^ input_b[1];
  assign cgp_core_073 = input_c[0] | input_h[0];
  assign cgp_core_075 = input_b[1] | cgp_core_066;
  assign cgp_core_076 = input_f[0] ^ input_i[1];
  assign cgp_core_077 = cgp_core_075 | cgp_core_071;
  assign cgp_core_078 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_079 = ~input_f[0];
  assign cgp_core_080_not = ~input_c[1];
  assign cgp_core_081 = ~(input_i[0] & input_d[0]);
  assign cgp_core_083 = ~input_e[1];
  assign cgp_core_084 = input_i[1] | input_g[1];
  assign cgp_core_085 = ~(input_f[0] & input_a[0]);
  assign cgp_core_086 = input_g[1] | input_g[0];
  assign cgp_core_088 = input_i[1] ^ input_g[0];
  assign cgp_core_089 = ~input_g[1];
  assign cgp_core_090 = input_h[0] & input_f[1];
  assign cgp_core_092 = ~cgp_core_077;
  assign cgp_core_093 = input_h[1] & cgp_core_092;
  assign cgp_core_094 = cgp_core_093 & input_i[1];
  assign cgp_core_095 = ~(input_c[1] | cgp_core_077);
  assign cgp_core_097 = input_e[1] | input_e[1];
  assign cgp_core_099 = input_d[1] & cgp_core_095;
  assign cgp_core_100 = ~(input_c[0] & input_f[1]);
  assign cgp_core_101 = input_a[1] ^ input_a[0];
  assign cgp_core_103 = ~(input_h[0] | input_c[0]);
  assign cgp_core_104 = ~(input_d[1] & input_d[1]);
  assign cgp_core_105 = input_e[0] | input_a[1];
  assign cgp_core_106 = ~(input_i[1] | input_f[1]);
  assign cgp_core_107 = cgp_core_099 | cgp_core_094;
  assign cgp_core_108 = ~(input_h[1] | input_g[1]);

  assign cgp_out[0] = cgp_core_107;
endmodule