module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018_not;
  wire cgp_core_019;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058_not;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069_not;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_018_not = ~input_e[2];
  assign cgp_core_019 = ~(input_e[1] & input_d[0]);
  assign cgp_core_022_not = ~input_b[2];
  assign cgp_core_023 = input_d[2] | input_d[0];
  assign cgp_core_024_not = ~input_c[1];
  assign cgp_core_026 = ~input_d[0];
  assign cgp_core_027 = ~input_e[0];
  assign cgp_core_028 = input_b[1] | input_a[1];
  assign cgp_core_030 = ~input_e[1];
  assign cgp_core_031 = ~(input_a[2] ^ input_a[1]);
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_034 = input_c[1] & input_b[1];
  assign cgp_core_035 = cgp_core_032 | cgp_core_034;
  assign cgp_core_038 = input_e[2] | cgp_core_035;
  assign cgp_core_039 = input_b[1] | input_c[1];
  assign cgp_core_042 = input_c[0] | input_e[2];
  assign cgp_core_045 = ~input_a[0];
  assign cgp_core_048 = ~(input_c[1] ^ input_c[1]);
  assign cgp_core_049 = input_a[2] & cgp_core_038;
  assign cgp_core_050_not = ~input_e[1];
  assign cgp_core_053 = ~(input_b[0] & input_a[2]);
  assign cgp_core_055 = input_c[2] | cgp_core_049;
  assign cgp_core_056 = input_e[1] & input_b[2];
  assign cgp_core_057 = input_b[2] | input_d[2];
  assign cgp_core_058_not = ~input_a[0];
  assign cgp_core_059 = ~cgp_core_057;
  assign cgp_core_060 = input_c[1] & input_b[2];
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_062 = cgp_core_061 & cgp_core_059;
  assign cgp_core_063 = ~(input_e[1] ^ input_b[1]);
  assign cgp_core_065 = input_a[2] & cgp_core_062;
  assign cgp_core_067 = input_d[2] ^ input_a[0];
  assign cgp_core_069_not = ~input_a[1];
  assign cgp_core_072 = ~(input_d[0] & input_c[2]);
  assign cgp_core_073 = ~(input_c[1] & input_b[2]);
  assign cgp_core_075 = ~(input_e[2] | input_e[0]);
  assign cgp_core_076 = ~(input_b[0] | input_b[1]);
  assign cgp_core_078 = input_c[1] | input_e[0];
  assign cgp_core_079 = input_d[2] | input_e[1];
  assign cgp_core_080 = input_c[1] & input_d[0];

  assign cgp_out[0] = cgp_core_065;
endmodule