module top #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 12,
parameter FEAT_BITS = 3,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1470


)(
    input   [FEAT_CNT * FEAT_BITS   -1:0] features,
    output  [$clog2(CLASS_CNT)      -1:0] prediction
);
localparam  SUM_BITS    = $clog2(HIDDEN_CNT + 1);
localparam  SCORE_BITS  = SUM_BITS + 1;
localparam  INDEX_BITS  = $clog2(FEAT_CNT + 1) + FEAT_BITS;

wire            [FEAT_BITS                  -1:0] feature_array [FEAT_CNT-1:0];
wire            [HIDDEN_CNT                 -1:0] hidden;
wire            [HIDDEN_CNT                 -1:0] hidden_n;
wire            [SUM_BITS                   -1:0] popcount      [CLASS_CNT-1:0]; 
wire            [(SUM_BITS + 1)             -1:0] scores        [CLASS_CNT-1:0]; 
wire            [CLASS_CNT * (SUM_BITS + 1) -1:0] score_vec; 

assign hidden_n = ~hidden;

genvar i;
generate
    for(i=0; i<FEAT_CNT; i=i+1) begin: l1
        assign feature_array[i] = features[i*FEAT_BITS +: FEAT_BITS];
    end
endgenerate
generate
    for(i=0;i<CLASS_CNT;i=i+1) begin: l2
        assign score_vec[i*SCORE_BITS +: SCORE_BITS] = scores[i];
    end
endgenerate



    ltg_0 ltg_0_hn (feature_array[3], feature_array[7], feature_array[10], hidden[0]);
    ltg_1 ltg_1_hn (feature_array[0], feature_array[2], feature_array[6], feature_array[7], feature_array[9], hidden[1]);
    ltg_2 ltg_2_hn (feature_array[0], feature_array[2], hidden[2]);
    ltg_3 ltg_3_hn (feature_array[1], feature_array[2], feature_array[3], feature_array[4], feature_array[9], feature_array[10], hidden[3]);
    ltg_4 ltg_4_hn (feature_array[0], feature_array[1], feature_array[2], feature_array[3], feature_array[8], hidden[4]);
    ltg_5 ltg_5_hn (feature_array[0], feature_array[2], feature_array[4], feature_array[5], feature_array[6], feature_array[9], hidden[5]);
assign hidden[6] = 1;
assign hidden[7] = 0;
    ltg_6 ltg_6_hn (feature_array[3], feature_array[6], feature_array[7], hidden[8]);
    ltg_7 ltg_7_hn (feature_array[2], feature_array[4], feature_array[8], feature_array[9], feature_array[10], hidden[9]);
assign hidden[10] = 0;
    ltg_8 ltg_8_hn (feature_array[1], feature_array[4], feature_array[7], feature_array[10], hidden[11]);
    
    popcount_0 popcount_0_pc ({hidden[11], hidden_n[10], hidden[9], hidden[8], hidden[7], hidden_n[6], hidden[5], hidden[4], hidden[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[0]);
    assign scores[0] = 2*popcount[0] + 0;

    popcount_1 popcount_1_pc ({hidden[11], hidden_n[10], hidden[9], hidden[8], hidden[7], hidden_n[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[1]);
    assign scores[1] = 2*popcount[1] + 0;

    popcount_2 popcount_2_pc ({hidden[11], hidden_n[10], hidden[9], hidden[8], hidden_n[7], hidden[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[2]);
    assign scores[2] = 2*popcount[2] + 0;

    popcount_3 popcount_3_pc ({hidden_n[11], hidden_n[10], hidden[9], hidden[8], hidden_n[7], hidden[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[3]);
    assign scores[3] = 2*popcount[3] + 0;

    popcount_4 popcount_4_pc ({hidden_n[11], hidden_n[10], hidden[9], hidden[8], hidden_n[7], hidden[6], hidden[5], hidden[4], hidden_n[3], hidden_n[2], hidden[1], hidden[0]}, popcount[4]);
    assign scores[4] = 2*popcount[4] + 0;

    popcount_5 popcount_5_pc ({hidden_n[11], hidden[10], hidden[9], hidden_n[8], hidden_n[7], hidden_n[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[5]);
    assign scores[5] = 2*popcount[5] + 0;

    popcount_6 popcount_6_pc ({hidden_n[11], hidden[10], hidden[9], hidden_n[8], hidden[7], hidden_n[6], hidden[5], hidden[4], hidden[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[6]);
    assign scores[6] = 2*popcount[6] + 0;



argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS+1)) result (
    .inx(score_vec),
    .outimax(prediction)
);
endmodule

module ltg_0(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_042;

  assign cgp_core_013 = input_a[0] & input_b[1];
  assign cgp_core_014 = input_b[1] & input_c[1];
  assign cgp_core_015 = input_b[1] ^ input_b[1];
  assign cgp_core_017 = cgp_core_014 | input_a[1];
  assign cgp_core_018 = input_a[2] | input_c[2];
  assign cgp_core_019 = input_a[2] & input_c[2];
  assign cgp_core_020 = cgp_core_018 | cgp_core_017;
  assign cgp_core_021 = cgp_core_018 & cgp_core_017;
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_023_not = ~input_a[1];
  assign cgp_core_024 = ~cgp_core_022;
  assign cgp_core_025 = ~cgp_core_020;
  assign cgp_core_026 = input_b[2] & cgp_core_025;
  assign cgp_core_028 = ~(input_b[2] ^ cgp_core_020);
  assign cgp_core_029 = cgp_core_028 & cgp_core_024;
  assign cgp_core_031 = input_c[2] | input_b[1];
  assign cgp_core_032 = input_b[1] & cgp_core_029;
  assign cgp_core_033 = ~(input_c[1] ^ input_a[1]);
  assign cgp_core_034 = input_a[1] & cgp_core_029;
  assign cgp_core_035 = ~input_b[0];
  assign cgp_core_037 = input_a[1] & cgp_core_034;
  assign cgp_core_040 = cgp_core_037 | cgp_core_032;
  assign cgp_core_042 = cgp_core_040 | cgp_core_026;

  assign cgp_out[0] = cgp_core_042;
endmodule
module ltg_1(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065_not;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_072_not;
  wire cgp_core_073;
  wire cgp_core_078;

  assign cgp_core_018 = input_e[0] ^ input_d[2];
  assign cgp_core_019 = input_e[0] | input_b[1];
  assign cgp_core_020 = ~(input_c[2] ^ input_b[2]);
  assign cgp_core_021 = ~(input_d[0] & input_c[1]);
  assign cgp_core_022 = ~input_b[0];
  assign cgp_core_023 = ~(input_a[0] ^ input_c[2]);
  assign cgp_core_024 = ~(input_d[2] & input_a[2]);
  assign cgp_core_025 = input_c[1] | input_e[0];
  assign cgp_core_026 = ~(input_b[1] & input_a[0]);
  assign cgp_core_028 = input_d[1] ^ input_a[0];
  assign cgp_core_029 = input_d[1] ^ input_e[1];
  assign cgp_core_030 = input_a[1] ^ input_c[1];
  assign cgp_core_032 = ~(input_a[0] ^ input_e[2]);
  assign cgp_core_033 = input_b[0] ^ input_a[2];
  assign cgp_core_035 = ~(input_e[2] | input_b[0]);
  assign cgp_core_037 = ~(input_b[0] | input_d[1]);
  assign cgp_core_039 = ~(input_d[1] ^ input_d[1]);
  assign cgp_core_041 = ~(input_b[2] | input_d[0]);
  assign cgp_core_042 = input_e[1] | input_b[0];
  assign cgp_core_043 = ~(input_b[1] & input_d[2]);
  assign cgp_core_044 = ~input_c[0];
  assign cgp_core_048 = ~(input_d[0] | input_c[2]);
  assign cgp_core_049 = input_e[1] ^ input_b[2];
  assign cgp_core_052 = input_c[2] ^ input_d[2];
  assign cgp_core_053 = ~(input_c[1] & input_d[2]);
  assign cgp_core_055 = ~input_e[1];
  assign cgp_core_058 = ~(input_c[2] | input_d[0]);
  assign cgp_core_060 = ~(input_d[1] & input_b[0]);
  assign cgp_core_061 = input_d[0] ^ input_a[0];
  assign cgp_core_063 = input_e[2] ^ input_b[2];
  assign cgp_core_064 = input_b[0] & input_c[1];
  assign cgp_core_065_not = ~input_a[2];
  assign cgp_core_066 = ~input_d[1];
  assign cgp_core_068 = ~input_a[0];
  assign cgp_core_069 = ~input_e[0];
  assign cgp_core_072_not = ~input_a[2];
  assign cgp_core_073 = ~(input_a[2] ^ input_e[0]);
  assign cgp_core_078 = ~(input_a[2] & input_c[0]);

  assign cgp_out[0] = cgp_core_024;
endmodule
module ltg_2(input [2:0] input_a, input [2:0] input_b, output [0:0] cgp_out);
  wire cgp_core_008;
  wire cgp_core_009;
  wire cgp_core_010;
  wire cgp_core_011;
  wire cgp_core_013;
  wire cgp_core_015_not;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_021;
  wire cgp_core_023;

  assign cgp_core_008 = ~input_b[2];
  assign cgp_core_009 = input_a[2] & cgp_core_008;
  assign cgp_core_010 = ~(input_a[2] ^ input_b[2]);
  assign cgp_core_011 = ~input_b[1];
  assign cgp_core_013 = cgp_core_011 & cgp_core_010;
  assign cgp_core_015_not = ~input_a[2];
  assign cgp_core_016 = ~(input_a[2] | input_b[2]);
  assign cgp_core_017 = input_a[0] & input_a[1];
  assign cgp_core_018 = cgp_core_017 & input_a[2];
  assign cgp_core_019_not = ~input_a[0];
  assign cgp_core_021 = cgp_core_018 | cgp_core_013;
  assign cgp_core_023 = cgp_core_021 | cgp_core_009;

  assign cgp_out[0] = cgp_core_023;
endmodule
module ltg_3(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088_not;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_098;

  assign cgp_core_020 = ~input_f[1];
  assign cgp_core_022 = input_a[1] ^ input_b[1];
  assign cgp_core_023 = input_a[1] & input_b[1];
  assign cgp_core_027 = input_a[2] ^ input_b[2];
  assign cgp_core_028 = input_a[2] & input_b[2];
  assign cgp_core_029 = cgp_core_027 ^ cgp_core_023;
  assign cgp_core_030 = cgp_core_027 & cgp_core_023;
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = ~(input_e[0] & input_f[0]);
  assign cgp_core_033 = ~(input_b[1] | input_d[0]);
  assign cgp_core_034 = input_c[1] ^ input_d[1];
  assign cgp_core_035 = input_a[1] | input_a[0];
  assign cgp_core_036 = ~cgp_core_034;
  assign cgp_core_037 = ~(input_f[2] | input_a[0]);
  assign cgp_core_038 = input_d[1] | input_c[1];
  assign cgp_core_039 = input_c[2] ^ input_d[2];
  assign cgp_core_040 = input_c[2] & input_d[2];
  assign cgp_core_041 = cgp_core_039 ^ cgp_core_038;
  assign cgp_core_042 = cgp_core_039 & cgp_core_038;
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;
  assign cgp_core_046 = input_e[1] | input_f[1];
  assign cgp_core_047 = input_e[1] & input_f[1];
  assign cgp_core_049 = ~(input_e[1] & input_c[0]);
  assign cgp_core_051 = input_e[2] | input_f[2];
  assign cgp_core_052 = input_a[0] & input_a[0];
  assign cgp_core_053 = cgp_core_051 | cgp_core_047;
  assign cgp_core_054 = ~(input_f[2] | input_f[1]);
  assign cgp_core_055 = ~(input_c[0] | input_c[1]);
  assign cgp_core_056 = input_f[2] | input_c[1];
  assign cgp_core_058 = cgp_core_036 ^ cgp_core_046;
  assign cgp_core_059 = cgp_core_036 & cgp_core_046;
  assign cgp_core_063 = cgp_core_041 ^ cgp_core_053;
  assign cgp_core_064 = cgp_core_041 & cgp_core_053;
  assign cgp_core_065 = cgp_core_063 ^ cgp_core_059;
  assign cgp_core_066 = cgp_core_063 & cgp_core_059;
  assign cgp_core_067 = cgp_core_064 | cgp_core_066;
  assign cgp_core_069 = input_f[2] & input_e[2];
  assign cgp_core_070 = cgp_core_043 | cgp_core_067;
  assign cgp_core_071 = cgp_core_043 & cgp_core_067;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;
  assign cgp_core_074 = ~cgp_core_072;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = cgp_core_031 & cgp_core_075;
  assign cgp_core_078 = ~(cgp_core_031 ^ cgp_core_070);
  assign cgp_core_079 = cgp_core_078 & cgp_core_074;
  assign cgp_core_080 = ~cgp_core_065;
  assign cgp_core_081 = cgp_core_029 & cgp_core_080;
  assign cgp_core_082 = cgp_core_081 & cgp_core_079;
  assign cgp_core_083 = ~(cgp_core_029 ^ cgp_core_065);
  assign cgp_core_084 = cgp_core_083 & cgp_core_079;
  assign cgp_core_085 = ~(input_f[0] ^ input_e[1]);
  assign cgp_core_087 = cgp_core_022 & cgp_core_084;
  assign cgp_core_088_not = ~cgp_core_058;
  assign cgp_core_089 = cgp_core_088_not & cgp_core_084;
  assign cgp_core_090 = input_b[2] | input_f[2];
  assign cgp_core_094 = input_c[0] & input_c[1];
  assign cgp_core_095 = cgp_core_087 | cgp_core_082;
  assign cgp_core_096 = cgp_core_089 | cgp_core_095;
  assign cgp_core_098 = cgp_core_096 | cgp_core_076;

  assign cgp_out[0] = cgp_core_098;
endmodule
module ltg_4(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_b[1] | input_c[0]);
  assign cgp_core_018 = ~(input_b[0] & input_d[0]);
  assign cgp_core_019 = ~input_e[0];
  assign cgp_core_024 = input_d[2] | input_d[2];
  assign cgp_core_026 = ~(input_c[0] & input_e[2]);
  assign cgp_core_027 = ~(input_a[1] ^ input_b[1]);
  assign cgp_core_028 = input_c[1] | input_a[1];
  assign cgp_core_029 = ~input_c[0];
  assign cgp_core_031 = input_e[2] | input_a[2];
  assign cgp_core_032 = input_d[1] & input_b[0];
  assign cgp_core_033 = input_b[0] | input_d[1];
  assign cgp_core_035 = ~input_a[1];
  assign cgp_core_036 = ~input_b[2];
  assign cgp_core_037 = input_d[2] ^ input_b[0];
  assign cgp_core_039 = input_d[1] ^ input_b[2];
  assign cgp_core_041 = ~input_d[2];
  assign cgp_core_045 = input_a[0] ^ input_c[2];
  assign cgp_core_048 = input_c[0] ^ input_b[1];
  assign cgp_core_049 = ~(cgp_core_026 & input_e[2]);
  assign cgp_core_050 = ~(input_e[2] | input_c[0]);
  assign cgp_core_051 = input_c[2] & input_b[1];
  assign cgp_core_055 = input_a[1] ^ input_d[1];
  assign cgp_core_057 = input_e[0] | input_a[0];
  assign cgp_core_058 = ~(input_a[2] & input_c[0]);
  assign cgp_core_059 = ~(input_d[2] & input_c[1]);
  assign cgp_core_061 = cgp_core_055 & input_e[0];
  assign cgp_core_062 = cgp_core_061 & input_d[2];
  assign cgp_core_063 = input_a[0] | input_c[1];
  assign cgp_core_064 = input_a[1] | input_a[2];
  assign cgp_core_066 = ~input_d[0];
  assign cgp_core_068 = ~(input_c[2] & cgp_core_045);
  assign cgp_core_069 = input_e[1] ^ input_b[1];
  assign cgp_core_070 = input_e[1] & input_d[2];
  assign cgp_core_072 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_073 = ~(input_d[1] ^ input_d[0]);
  assign cgp_core_075 = ~(input_e[0] & cgp_core_072);
  assign cgp_core_076 = ~input_c[1];
  assign cgp_core_079 = input_c[1] ^ input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule
module ltg_5(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_020 = input_c[0] ^ input_e[0];
  assign cgp_core_021 = input_c[0] & input_e[0];
  assign cgp_core_023 = input_c[1] & input_e[1];
  assign cgp_core_027 = input_c[2] ^ input_e[2];
  assign cgp_core_028 = input_c[2] & input_b[0];
  assign cgp_core_029 = ~input_f[0];
  assign cgp_core_030 = input_f[2] & cgp_core_023;
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = input_a[0] ^ cgp_core_020;
  assign cgp_core_033 = input_a[0] & cgp_core_020;
  assign cgp_core_034 = input_a[1] ^ cgp_core_021;
  assign cgp_core_035 = input_a[1] & cgp_core_021;
  assign cgp_core_036 = cgp_core_034 ^ input_b[0];
  assign cgp_core_037 = cgp_core_034 & input_d[2];
  assign cgp_core_038 = cgp_core_035 | cgp_core_037;
  assign cgp_core_039 = input_a[2] ^ cgp_core_029;
  assign cgp_core_040 = input_a[2] & cgp_core_029;
  assign cgp_core_041 = cgp_core_039 ^ cgp_core_038;
  assign cgp_core_042 = cgp_core_039 & cgp_core_038;
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;
  assign cgp_core_044 = cgp_core_031 ^ cgp_core_043;
  assign cgp_core_045 = cgp_core_031 & cgp_core_043;
  assign cgp_core_047 = input_d[0] & input_f[0];
  assign cgp_core_048 = input_d[1] ^ input_f[1];
  assign cgp_core_049 = input_d[1] & input_f[1];
  assign cgp_core_050 = cgp_core_048 ^ cgp_core_047;
  assign cgp_core_051 = cgp_core_048 & cgp_core_047;
  assign cgp_core_052 = cgp_core_049 | cgp_core_051;
  assign cgp_core_053 = input_d[2] ^ input_f[2];
  assign cgp_core_054 = input_d[2] & input_f[2];
  assign cgp_core_055 = cgp_core_053 ^ cgp_core_052;
  assign cgp_core_056 = cgp_core_053 & cgp_core_052;
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058 = input_b[0] ^ input_b[1];
  assign cgp_core_059 = input_b[0] & input_b[1];
  assign cgp_core_060 = ~(input_b[1] & cgp_core_050);
  assign cgp_core_061 = input_b[1] & cgp_core_050;
  assign cgp_core_062 = ~(cgp_core_060 & cgp_core_059);
  assign cgp_core_063 = cgp_core_060 & cgp_core_059;
  assign cgp_core_064 = input_f[1] | cgp_core_063;
  assign cgp_core_065 = input_b[2] ^ cgp_core_055;
  assign cgp_core_066 = input_b[2] & cgp_core_055;
  assign cgp_core_067 = cgp_core_065 ^ input_d[0];
  assign cgp_core_068 = cgp_core_065 & cgp_core_064;
  assign cgp_core_069 = cgp_core_066 | cgp_core_068;
  assign cgp_core_070 = cgp_core_057 ^ cgp_core_069;
  assign cgp_core_071 = cgp_core_057 & cgp_core_069;
  assign cgp_core_072 = ~cgp_core_071;
  assign cgp_core_073 = cgp_core_045 & cgp_core_072;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = cgp_core_044 & cgp_core_075;
  assign cgp_core_078 = ~(cgp_core_044 ^ cgp_core_070);
  assign cgp_core_080 = ~cgp_core_067;
  assign cgp_core_081 = cgp_core_041 & cgp_core_080;
  assign cgp_core_082 = cgp_core_081 & cgp_core_078;
  assign cgp_core_083 = cgp_core_041 & cgp_core_067;
  assign cgp_core_084 = cgp_core_083 & cgp_core_078;
  assign cgp_core_085 = ~cgp_core_062;
  assign cgp_core_086 = cgp_core_036 & cgp_core_085;
  assign cgp_core_087 = cgp_core_086 & cgp_core_084;
  assign cgp_core_088 = cgp_core_036 & cgp_core_062;
  assign cgp_core_089 = cgp_core_088 & cgp_core_084;
  assign cgp_core_090 = ~cgp_core_058;
  assign cgp_core_091 = cgp_core_032 & cgp_core_090;
  assign cgp_core_092 = input_c[1] & cgp_core_089;
  assign cgp_core_093 = ~(cgp_core_032 ^ cgp_core_058);
  assign cgp_core_094 = input_d[1] & cgp_core_089;
  assign cgp_core_095 = cgp_core_087 | cgp_core_082;
  assign cgp_core_096 = cgp_core_092 | cgp_core_095;
  assign cgp_core_097 = cgp_core_073 | cgp_core_094;
  assign cgp_core_098 = cgp_core_076 | cgp_core_097;
  assign cgp_core_099 = cgp_core_096 | cgp_core_098;

  assign cgp_out[0] = input_e[2];
endmodule
module ltg_6(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;

  assign cgp_core_011 = input_a[0] ^ input_b[0];
  assign cgp_core_012 = input_a[0] & input_b[0];
  assign cgp_core_013 = input_a[1] ^ input_b[1];
  assign cgp_core_014 = input_a[1] & input_b[1];
  assign cgp_core_015 = cgp_core_013 ^ cgp_core_012;
  assign cgp_core_016 = cgp_core_013 & cgp_core_012;
  assign cgp_core_017 = ~(cgp_core_014 | cgp_core_016);
  assign cgp_core_018 = input_a[2] ^ input_b[2];
  assign cgp_core_019 = input_a[2] & input_b[2];
  assign cgp_core_020 = ~(cgp_core_018 & cgp_core_017);
  assign cgp_core_021 = cgp_core_018 & cgp_core_017;
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_023 = ~cgp_core_022;
  assign cgp_core_024 = ~input_c[2];
  assign cgp_core_025 = cgp_core_020 & cgp_core_024;
  assign cgp_core_026 = cgp_core_025 & cgp_core_023;
  assign cgp_core_027 = ~(cgp_core_020 ^ input_c[2]);
  assign cgp_core_028 = cgp_core_027 & cgp_core_023;
  assign cgp_core_029 = ~input_c[1];
  assign cgp_core_032 = ~cgp_core_015;
  assign cgp_core_033 = cgp_core_032 & cgp_core_028;
  assign cgp_core_034 = ~input_c[0];
  assign cgp_core_035 = cgp_core_011 & cgp_core_034;
  assign cgp_core_036 = cgp_core_035 & cgp_core_033;
  assign cgp_core_037 = ~(input_c[0] ^ input_c[0]);
  assign cgp_core_038 = cgp_core_037 & cgp_core_033;
  assign cgp_core_040 = cgp_core_022 | cgp_core_038;
  assign cgp_core_041 = cgp_core_026 | cgp_core_040;

  assign cgp_out[0] = 1'b1;
endmodule
module ltg_7(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_a[2] & input_a[2]);
  assign cgp_core_019 = ~input_b[1];
  assign cgp_core_024 = input_c[2] | input_d[2];
  assign cgp_core_026 = input_e[0] ^ input_b[0];
  assign cgp_core_027 = ~input_b[0];
  assign cgp_core_028 = ~input_c[1];
  assign cgp_core_030 = ~(input_c[1] | input_b[0]);
  assign cgp_core_034 = ~(input_e[1] & input_b[1]);
  assign cgp_core_036 = ~(input_c[0] & input_c[2]);
  assign cgp_core_038 = ~input_c[2];
  assign cgp_core_040 = input_e[0] & input_d[1];
  assign cgp_core_041 = input_e[2] ^ input_b[2];
  assign cgp_core_042 = ~input_c[2];
  assign cgp_core_044 = input_d[2] | input_e[1];
  assign cgp_core_046_not = ~input_b[1];
  assign cgp_core_049 = ~(input_c[2] | input_e[2]);
  assign cgp_core_050 = ~(input_a[1] | input_e[1]);
  assign cgp_core_051 = input_c[0] & input_d[1];
  assign cgp_core_058 = input_e[2] | input_b[0];
  assign cgp_core_059 = ~input_b[1];
  assign cgp_core_060 = input_a[2] & input_b[1];
  assign cgp_core_061 = ~(input_b[1] | input_b[1]);
  assign cgp_core_063 = ~(input_d[2] | input_d[2]);
  assign cgp_core_064 = ~(input_e[1] & input_c[2]);
  assign cgp_core_065 = ~(input_a[2] | input_a[2]);
  assign cgp_core_067 = ~(input_c[2] | input_d[0]);
  assign cgp_core_068 = ~input_e[1];
  assign cgp_core_070 = ~(input_d[2] & input_e[1]);
  assign cgp_core_072 = ~(input_b[2] & input_b[2]);
  assign cgp_core_076 = ~input_d[0];
  assign cgp_core_078 = ~(input_d[1] ^ input_c[0]);
  assign cgp_core_079 = input_c[1] ^ input_c[2];

  assign cgp_out[0] = cgp_core_049;
endmodule
module ltg_8(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_015 = input_c[2] ^ input_d[0];
  assign cgp_core_016 = ~input_b[2];
  assign cgp_core_019 = ~input_c[0];
  assign cgp_core_020 = input_a[1] | input_b[1];
  assign cgp_core_021 = input_a[2] ^ input_b[2];
  assign cgp_core_022 = input_a[2] & input_b[2];
  assign cgp_core_023 = cgp_core_021 ^ cgp_core_020;
  assign cgp_core_024 = cgp_core_021 & cgp_core_020;
  assign cgp_core_025 = cgp_core_022 | cgp_core_024;
  assign cgp_core_026 = input_d[2] & input_b[0];
  assign cgp_core_027 = ~input_d[0];
  assign cgp_core_028 = ~(input_d[2] & input_b[0]);
  assign cgp_core_029 = input_c[1] & input_d[1];
  assign cgp_core_030 = input_c[0] & input_d[0];
  assign cgp_core_033 = input_c[2] ^ input_d[2];
  assign cgp_core_034 = input_c[2] & input_d[2];
  assign cgp_core_035 = cgp_core_033 ^ cgp_core_029;
  assign cgp_core_036 = cgp_core_033 & cgp_core_029;
  assign cgp_core_037 = cgp_core_034 | cgp_core_036;
  assign cgp_core_038 = ~cgp_core_037;
  assign cgp_core_039 = cgp_core_025 & cgp_core_038;
  assign cgp_core_040 = ~(cgp_core_025 ^ cgp_core_037);
  assign cgp_core_041 = ~cgp_core_035;
  assign cgp_core_042 = cgp_core_023 & cgp_core_041;
  assign cgp_core_043 = cgp_core_042 & cgp_core_040;
  assign cgp_core_045 = ~input_d[2];
  assign cgp_core_046 = input_a[1] | input_c[0];
  assign cgp_core_048 = ~(input_c[1] ^ input_d[0]);
  assign cgp_core_050_not = ~input_c[2];
  assign cgp_core_051 = ~(input_b[0] ^ input_b[0]);
  assign cgp_core_052 = ~(input_b[1] ^ input_d[1]);
  assign cgp_core_053_not = ~input_b[1];
  assign cgp_core_054 = ~input_c[2];
  assign cgp_core_058 = cgp_core_043 | cgp_core_039;
  assign cgp_core_059 = ~(input_c[0] ^ input_d[2]);

  assign cgp_out[0] = cgp_core_058;
endmodule
module popcount_0(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067_not;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~(input_a[8] | input_a[9]);
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_025 = input_a[6] ^ input_a[0];
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[7] | input_a[9]);
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_043 = ~(input_a[9] & input_a[1]);
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_049 = ~input_a[8];
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 | cgp_core_063;
  assign cgp_core_067_not = ~input_a[9];
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_065;
  assign cgp_core_072 = cgp_core_069 & cgp_core_065;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~(input_a[10] & input_a[7]);
  assign cgp_core_075 = input_a[0] | input_a[9];
  assign cgp_core_077 = ~input_a[9];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_1(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035_not;
  wire cgp_core_038_not;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = ~(input_a[1] & input_a[3]);
  assign cgp_core_015 = ~(input_a[1] | input_a[1]);
  assign cgp_core_016 = ~input_a[7];
  assign cgp_core_019 = ~input_a[3];
  assign cgp_core_020 = input_a[11] ^ input_a[6];
  assign cgp_core_023 = ~(input_a[3] ^ input_a[5]);
  assign cgp_core_024 = ~input_a[3];
  assign cgp_core_026 = ~(input_a[9] & input_a[1]);
  assign cgp_core_027 = ~(input_a[11] ^ input_a[10]);
  assign cgp_core_028 = ~(input_a[11] | input_a[6]);
  assign cgp_core_031 = input_a[1] ^ input_a[11];
  assign cgp_core_032 = ~input_a[4];
  assign cgp_core_033 = ~(input_a[6] & input_a[10]);
  assign cgp_core_035_not = ~input_a[3];
  assign cgp_core_038_not = ~input_a[1];
  assign cgp_core_041 = ~(input_a[0] ^ input_a[8]);
  assign cgp_core_042 = ~(input_a[4] & input_a[9]);
  assign cgp_core_045 = ~(input_a[3] ^ input_a[7]);
  assign cgp_core_046 = input_a[1] & input_a[10];
  assign cgp_core_049 = ~(input_a[11] | input_a[9]);
  assign cgp_core_051 = input_a[7] | input_a[2];
  assign cgp_core_052 = ~(input_a[1] & input_a[5]);
  assign cgp_core_053 = ~(input_a[2] ^ input_a[8]);
  assign cgp_core_054 = ~(input_a[1] | input_a[2]);
  assign cgp_core_057 = ~(input_a[7] & input_a[0]);
  assign cgp_core_061 = ~input_a[0];
  assign cgp_core_063 = ~(input_a[8] ^ input_a[4]);
  assign cgp_core_065 = input_a[1] | input_a[6];
  assign cgp_core_066 = ~input_a[3];
  assign cgp_core_067 = ~(input_a[0] & input_a[6]);
  assign cgp_core_068 = ~input_a[10];
  assign cgp_core_069 = ~(input_a[7] ^ input_a[3]);
  assign cgp_core_071 = ~(input_a[4] | input_a[9]);
  assign cgp_core_072 = ~input_a[7];
  assign cgp_core_075 = input_a[2] ^ input_a[5];
  assign cgp_core_077 = ~(input_a[3] | input_a[8]);
  assign cgp_core_078 = input_a[9] ^ input_a[4];

  assign cgp_out[0] = 1'b0;
  assign cgp_out[1] = 1'b1;
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = 1'b0;
endmodule
module popcount_2(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_3(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055_not;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[9];
  assign cgp_core_020 = input_a[4] | input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = ~(input_a[2] & input_a[3]);
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_025 = ~(input_a[5] | input_a[2]);
  assign cgp_core_026 = ~cgp_core_016;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_016;
  assign cgp_core_031 = cgp_core_028 & cgp_core_016;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[7] | input_a[2]);
  assign cgp_core_036_not = ~input_a[2];
  assign cgp_core_038 = ~input_a[4];
  assign cgp_core_039 = input_a[1] ^ input_a[11];
  assign cgp_core_040 = ~(input_a[2] & input_a[5]);
  assign cgp_core_042 = input_a[7] & input_a[8];
  assign cgp_core_043 = ~(input_a[2] | input_a[2]);
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_047 = input_a[9] & input_a[6];
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_049 = ~input_a[7];
  assign cgp_core_050 = input_a[10] | input_a[9];
  assign cgp_core_051 = ~(input_a[3] | input_a[5]);
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_055_not = ~input_a[9];
  assign cgp_core_058 = ~(input_a[9] | input_a[6]);
  assign cgp_core_061 = input_a[4] ^ input_a[5];
  assign cgp_core_062 = input_a[1] | input_a[3];
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_052;
  assign cgp_core_065 = cgp_core_030 & cgp_core_052;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_026;
  assign cgp_core_067 = cgp_core_064 & cgp_core_026;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_053;
  assign cgp_core_070 = cgp_core_032 & cgp_core_053;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~(input_a[10] | input_a[7]);
  assign cgp_core_076 = input_a[8] ^ input_a[3];
  assign cgp_core_078 = input_a[1] | input_a[9];

  assign cgp_out[0] = cgp_core_016;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_4(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021_not;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_037_not;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_017_not = ~input_a[6];
  assign cgp_core_018 = input_a[2] ^ input_a[1];
  assign cgp_core_019 = input_a[5] ^ input_a[8];
  assign cgp_core_021_not = ~input_a[0];
  assign cgp_core_025 = input_a[1] & input_a[9];
  assign cgp_core_028 = input_a[8] & input_a[11];
  assign cgp_core_030 = ~(input_a[5] & input_a[3]);
  assign cgp_core_031 = input_a[3] & input_a[5];
  assign cgp_core_034 = input_a[11] | input_a[11];
  assign cgp_core_037_not = ~input_a[10];
  assign cgp_core_039 = ~(input_a[3] | input_a[11]);
  assign cgp_core_041 = input_a[1] | input_a[1];
  assign cgp_core_042 = input_a[6] | input_a[0];
  assign cgp_core_045 = input_a[11] & input_a[9];
  assign cgp_core_046 = ~(input_a[8] & input_a[1]);
  assign cgp_core_047 = input_a[10] & input_a[1];
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_049_not = ~input_a[11];
  assign cgp_core_051 = ~(input_a[8] ^ input_a[9]);
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_058 = input_a[8] & input_a[2];
  assign cgp_core_061 = ~input_a[2];
  assign cgp_core_063 = input_a[7] & input_a[8];
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_052;
  assign cgp_core_065 = cgp_core_030 & cgp_core_052;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_031 ^ cgp_core_053;
  assign cgp_core_070 = cgp_core_031 & cgp_core_053;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[11];
  assign cgp_core_075 = input_a[0] ^ input_a[3];
  assign cgp_core_076 = ~(input_a[3] & input_a[3]);
  assign cgp_core_077 = ~input_a[3];
  assign cgp_core_078 = ~(input_a[1] ^ input_a[11]);

  assign cgp_out[0] = input_a[4];
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_5(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_025 = input_a[11] & input_a[7];
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_037 = input_a[8] | input_a[3];
  assign cgp_core_038 = input_a[7] | input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[0] | input_a[3];
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] | input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = ~(input_a[9] | input_a[7]);
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_062 = ~cgp_core_026;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_052;
  assign cgp_core_065 = cgp_core_030 & cgp_core_052;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_026;
  assign cgp_core_067 = cgp_core_064 & cgp_core_026;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_053;
  assign cgp_core_070 = cgp_core_032 & cgp_core_053;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_076 = ~(input_a[9] ^ input_a[0]);
  assign cgp_core_077 = input_a[0] & input_a[8];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_6(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021_not;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_037_not;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_017_not = ~input_a[6];
  assign cgp_core_018 = input_a[2] ^ input_a[1];
  assign cgp_core_019 = input_a[5] ^ input_a[8];
  assign cgp_core_021_not = ~input_a[0];
  assign cgp_core_025 = input_a[1] & input_a[9];
  assign cgp_core_028 = input_a[8] & input_a[11];
  assign cgp_core_030 = ~(input_a[5] & input_a[3]);
  assign cgp_core_031 = input_a[3] & input_a[5];
  assign cgp_core_034 = input_a[11] | input_a[11];
  assign cgp_core_037_not = ~input_a[10];
  assign cgp_core_039 = ~(input_a[3] | input_a[11]);
  assign cgp_core_041 = input_a[1] | input_a[1];
  assign cgp_core_042 = input_a[6] | input_a[0];
  assign cgp_core_045 = input_a[11] & input_a[9];
  assign cgp_core_046 = ~(input_a[8] & input_a[1]);
  assign cgp_core_047 = input_a[10] & input_a[1];
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_049_not = ~input_a[11];
  assign cgp_core_051 = ~(input_a[8] ^ input_a[9]);
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_058 = input_a[8] & input_a[2];
  assign cgp_core_061 = ~input_a[2];
  assign cgp_core_063 = input_a[7] & input_a[8];
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_052;
  assign cgp_core_065 = cgp_core_030 & cgp_core_052;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_031 ^ cgp_core_053;
  assign cgp_core_070 = cgp_core_031 & cgp_core_053;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[11];
  assign cgp_core_075 = input_a[0] ^ input_a[3];
  assign cgp_core_076 = ~(input_a[3] & input_a[3]);
  assign cgp_core_077 = ~input_a[3];
  assign cgp_core_078 = ~(input_a[1] ^ input_a[11]);

  assign cgp_out[0] = input_a[4];
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module argmax #(
    parameter SIZE = 9,
    parameter BITS = 4,
    parameter INDEX_BITS = 4
) (
    input [SIZE*BITS-1:0] inx,
    output [INDEX_BITS-1:0] outimax
);

wire [INDEX_BITS-1:0] interm_argmax [SIZE-1:0];
wire [BITS-1:0] interm_max [SIZE-1:0];

assign interm_max[0] = inx[0+:BITS];
assign interm_argmax[0] = 0;

genvar j;
generate
for (j = 1; j < SIZE; j = j + 1) begin : whatss
	wire huge; //Flag that tracks if current sample is largest so far
	assign huge = inx[j*BITS+:BITS] > interm_max[j-1];
	assign interm_max[j] = huge ? inx[j*BITS+:BITS]:interm_max[j-1]; 
	assign interm_argmax[j] = huge ? j:interm_argmax[j-1];
end
endgenerate

assign outimax = interm_argmax[SIZE-1];

endmodule
