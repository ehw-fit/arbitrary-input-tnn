module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;

  assign cgp_core_016 = input_c[1] & input_e[0];
  assign cgp_core_017 = input_c[0] & input_f[1];
  assign cgp_core_018 = input_a[0] ^ input_g[0];
  assign cgp_core_022 = input_e[0] | input_c[0];
  assign cgp_core_023 = input_a[0] & input_f[1];
  assign cgp_core_024 = input_c[1] ^ cgp_core_016;
  assign cgp_core_027 = input_g[0] ^ cgp_core_024;
  assign cgp_core_028 = input_g[0] ^ input_e[1];
  assign cgp_core_030 = input_a[0] | input_a[1];
  assign cgp_core_031 = ~(input_b[1] & input_d[0]);
  assign cgp_core_032 = input_a[1] ^ input_d[0];
  assign cgp_core_033 = ~input_a[1];
  assign cgp_core_035 = ~(input_b[1] ^ input_d[1]);
  assign cgp_core_036 = ~(input_d[1] ^ cgp_core_033);
  assign cgp_core_037 = input_d[1] & cgp_core_033;
  assign cgp_core_038 = input_c[0] ^ input_f[0];
  assign cgp_core_039 = ~(input_e[0] & input_g[1]);
  assign cgp_core_041_not = ~input_f[0];
  assign cgp_core_042 = ~(input_f[1] ^ input_d[0]);
  assign cgp_core_043 = input_b[0] ^ input_g[0];
  assign cgp_core_045 = input_f[0] | input_g[1];
  assign cgp_core_047 = cgp_core_032 & input_c[0];
  assign cgp_core_049 = ~(input_a[0] | cgp_core_043);
  assign cgp_core_050_not = ~input_d[1];
  assign cgp_core_051 = ~input_g[1];
  assign cgp_core_052 = input_d[1] | input_g[0];
  assign cgp_core_053 = input_b[0] ^ input_b[1];
  assign cgp_core_056 = cgp_core_053 & input_a[1];
  assign cgp_core_058 = ~input_g[1];
  assign cgp_core_059 = ~(input_d[0] & input_g[1]);
  assign cgp_core_060 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_061 = ~input_e[0];
  assign cgp_core_062 = ~(input_c[1] & cgp_core_061);
  assign cgp_core_063 = cgp_core_062 & cgp_core_060;
  assign cgp_core_065 = ~(input_c[1] & cgp_core_060);
  assign cgp_core_066 = input_f[1] ^ input_c[1];
  assign cgp_core_070 = input_f[0] & input_d[0];
  assign cgp_core_072 = cgp_core_023 & input_g[1];
  assign cgp_core_073 = input_e[1] ^ cgp_core_070;
  assign cgp_core_074 = ~(cgp_core_023 ^ cgp_core_039);
  assign cgp_core_075 = input_c[0] | cgp_core_070;
  assign cgp_core_077 = cgp_core_059 | cgp_core_075;

  assign cgp_out[0] = 1'b0;
endmodule