module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051_not;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_077;

  assign cgp_core_015 = ~(input_a[6] & input_a[6]);
  assign cgp_core_016 = ~(input_a[7] | input_a[2]);
  assign cgp_core_017 = ~input_a[0];
  assign cgp_core_020 = input_a[11] | input_a[6];
  assign cgp_core_022 = input_a[5] & input_a[9];
  assign cgp_core_024 = ~(input_a[9] & input_a[0]);
  assign cgp_core_026 = ~input_a[10];
  assign cgp_core_027 = ~(input_a[9] | input_a[7]);
  assign cgp_core_028 = input_a[0] | input_a[10];
  assign cgp_core_030 = ~input_a[3];
  assign cgp_core_031 = input_a[3] ^ input_a[11];
  assign cgp_core_034 = input_a[1] ^ input_a[7];
  assign cgp_core_035 = input_a[6] & input_a[4];
  assign cgp_core_037 = ~input_a[7];
  assign cgp_core_038 = ~(input_a[0] | input_a[0]);
  assign cgp_core_040 = input_a[7] ^ input_a[8];
  assign cgp_core_042 = input_a[8] & input_a[10];
  assign cgp_core_044 = input_a[5] & input_a[10];
  assign cgp_core_046 = ~(input_a[7] & input_a[0]);
  assign cgp_core_047 = ~input_a[11];
  assign cgp_core_048 = input_a[1] | input_a[6];
  assign cgp_core_050 = input_a[11] & input_a[6];
  assign cgp_core_051_not = ~input_a[8];
  assign cgp_core_052 = ~(cgp_core_042 & cgp_core_048);
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_063 = ~(input_a[10] ^ input_a[1]);
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_052;
  assign cgp_core_065 = input_a[0] & input_a[6];
  assign cgp_core_069 = ~(input_a[3] & cgp_core_053);
  assign cgp_core_070 = input_a[3] & cgp_core_053;
  assign cgp_core_071 = ~(input_a[5] | input_a[7]);
  assign cgp_core_073 = input_a[2] | input_a[2];
  assign cgp_core_074 = input_a[2] & input_a[11];
  assign cgp_core_077 = input_a[2] & input_a[4];

  assign cgp_out[0] = input_a[7];
  assign cgp_out[1] = cgp_core_064;
  assign cgp_out[2] = cgp_core_069;
  assign cgp_out[3] = cgp_core_070;
endmodule