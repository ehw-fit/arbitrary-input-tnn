module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_036_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068_not;
  wire cgp_core_070;

  assign cgp_core_016 = input_b[1] | input_b[0];
  assign cgp_core_018 = ~(input_a[0] ^ input_e[1]);
  assign cgp_core_021 = input_b[1] | input_f[0];
  assign cgp_core_023 = ~(input_d[1] & input_b[0]);
  assign cgp_core_024 = ~(input_a[1] | input_b[1]);
  assign cgp_core_025_not = ~input_f[1];
  assign cgp_core_026 = ~input_a[0];
  assign cgp_core_027_not = ~input_f[1];
  assign cgp_core_030 = input_b[1] & input_c[0];
  assign cgp_core_032 = ~input_d[1];
  assign cgp_core_036_not = ~input_a[0];
  assign cgp_core_037 = input_c[0] | input_c[1];
  assign cgp_core_038 = input_e[1] & input_d[0];
  assign cgp_core_039 = ~(input_e[0] ^ input_b[0]);
  assign cgp_core_040 = ~(input_b[1] | input_e[0]);
  assign cgp_core_041 = input_f[1] ^ input_a[1];
  assign cgp_core_042 = ~(input_c[0] ^ input_f[0]);
  assign cgp_core_045 = ~(input_e[0] & input_d[0]);
  assign cgp_core_046 = input_e[1] & input_d[1];
  assign cgp_core_047 = ~input_e[1];
  assign cgp_core_051 = ~input_f[0];
  assign cgp_core_053 = ~(input_e[0] ^ input_d[0]);
  assign cgp_core_054 = input_c[0] | input_e[0];
  assign cgp_core_056 = input_e[1] | input_f[1];
  assign cgp_core_059 = ~(input_d[0] | input_c[1]);
  assign cgp_core_060 = ~(input_c[0] & input_e[0]);
  assign cgp_core_061 = input_b[0] | input_b[1];
  assign cgp_core_064 = ~(input_c[1] ^ input_a[1]);
  assign cgp_core_066 = ~(input_b[0] & input_a[0]);
  assign cgp_core_068_not = ~input_b[0];
  assign cgp_core_070 = input_c[1] ^ input_a[0];

  assign cgp_out[0] = 1'b1;
endmodule