module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055_not;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = input_b[0] | input_e[0];
  assign cgp_core_018 = input_b[0] & input_c[0];
  assign cgp_core_019 = input_b[1] ^ input_c[1];
  assign cgp_core_020 = input_b[1] & input_c[1];
  assign cgp_core_022 = cgp_core_019 & cgp_core_018;
  assign cgp_core_024 = input_b[2] ^ input_c[2];
  assign cgp_core_025 = input_c[1] & input_c[2];
  assign cgp_core_026 = input_a[2] ^ input_d[0];
  assign cgp_core_027 = cgp_core_024 & input_d[0];
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_029 = input_d[0] ^ input_e[0];
  assign cgp_core_030 = input_d[0] ^ input_e[0];
  assign cgp_core_031 = input_d[1] ^ input_e[1];
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_033 = cgp_core_031 ^ cgp_core_030;
  assign cgp_core_036 = input_d[2] ^ input_e[2];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_039 = cgp_core_036 & cgp_core_032;
  assign cgp_core_040 = cgp_core_037 | input_d[1];
  assign cgp_core_041 = cgp_core_017 ^ input_b[0];
  assign cgp_core_044 = ~(cgp_core_018 & cgp_core_033);
  assign cgp_core_047 = input_b[0] | input_e[2];
  assign cgp_core_048 = cgp_core_026 ^ cgp_core_036;
  assign cgp_core_049 = input_d[2] & cgp_core_036;
  assign cgp_core_050 = cgp_core_048 ^ input_c[0];
  assign cgp_core_052 = cgp_core_049 | input_a[1];
  assign cgp_core_054 = cgp_core_028 & cgp_core_040;
  assign cgp_core_055_not = ~cgp_core_052;
  assign cgp_core_057 = input_b[2] | cgp_core_052;
  assign cgp_core_058 = ~input_d[2];
  assign cgp_core_059 = ~cgp_core_057;
  assign cgp_core_060 = ~cgp_core_055_not;
  assign cgp_core_061 = ~cgp_core_055_not;
  assign cgp_core_062 = cgp_core_061 & cgp_core_059;
  assign cgp_core_063 = ~cgp_core_050;
  assign cgp_core_064 = input_a[2] & input_d[2];
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066 = input_a[2] ^ cgp_core_050;
  assign cgp_core_070 = input_a[1] & cgp_core_062;
  assign cgp_core_072 = input_a[1] & cgp_core_062;
  assign cgp_core_073 = ~cgp_core_041;
  assign cgp_core_074 = ~(input_a[0] | cgp_core_073);
  assign cgp_core_075 = cgp_core_074 & cgp_core_072;
  assign cgp_core_078 = cgp_core_070 | cgp_core_065;
  assign cgp_core_079 = cgp_core_075 | cgp_core_078;

  assign cgp_out[0] = 1'b0;
endmodule