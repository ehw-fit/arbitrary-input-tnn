module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052_not;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062_not;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_078_not;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_018 = ~input_a[2];
  assign cgp_core_019 = ~(input_d[1] ^ input_d[2]);
  assign cgp_core_020 = ~input_b[1];
  assign cgp_core_021 = ~(input_e[2] ^ input_a[0]);
  assign cgp_core_024 = ~(input_e[1] | input_e[1]);
  assign cgp_core_025 = ~(input_c[2] & input_a[2]);
  assign cgp_core_026 = ~input_d[0];
  assign cgp_core_027 = ~(input_e[0] & input_a[2]);
  assign cgp_core_028 = input_b[1] ^ input_e[2];
  assign cgp_core_030 = input_e[0] | input_c[0];
  assign cgp_core_033 = ~(input_e[2] & input_d[0]);
  assign cgp_core_034 = ~input_a[1];
  assign cgp_core_035 = ~input_c[1];
  assign cgp_core_036 = input_a[2] | input_a[1];
  assign cgp_core_039 = input_a[1] | input_e[0];
  assign cgp_core_041 = ~input_c[0];
  assign cgp_core_042 = ~input_c[2];
  assign cgp_core_043 = ~input_d[2];
  assign cgp_core_045 = ~(input_c[2] & input_e[2]);
  assign cgp_core_046 = input_b[2] ^ input_b[1];
  assign cgp_core_047 = ~(input_c[1] | input_c[1]);
  assign cgp_core_048 = input_e[2] ^ input_e[2];
  assign cgp_core_050 = ~input_a[1];
  assign cgp_core_052_not = ~input_d[1];
  assign cgp_core_053 = ~input_d[0];
  assign cgp_core_055 = input_b[0] ^ input_d[1];
  assign cgp_core_056 = input_b[1] ^ input_a[1];
  assign cgp_core_057 = ~(input_e[0] ^ input_e[2]);
  assign cgp_core_059 = input_d[0] ^ input_b[1];
  assign cgp_core_061 = input_c[1] & input_e[0];
  assign cgp_core_062_not = ~input_a[2];
  assign cgp_core_063 = input_b[1] & input_b[2];
  assign cgp_core_064 = cgp_core_063 & input_a[2];
  assign cgp_core_066 = ~(input_c[0] ^ input_d[0]);
  assign cgp_core_069 = ~(input_b[0] ^ input_c[1]);
  assign cgp_core_071 = ~(input_e[2] & input_b[2]);
  assign cgp_core_073 = ~(input_b[0] & input_b[2]);
  assign cgp_core_074 = ~(input_a[2] | input_d[2]);
  assign cgp_core_076 = ~(input_d[1] ^ input_c[0]);
  assign cgp_core_078_not = ~input_c[0];
  assign cgp_core_079 = ~(input_d[0] | input_e[2]);
  assign cgp_core_080 = input_c[1] & input_d[1];

  assign cgp_out[0] = cgp_core_064;
endmodule