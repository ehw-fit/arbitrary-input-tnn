module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_046_not;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052_not;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_088;
  wire cgp_core_091;
  wire cgp_core_094;
  wire cgp_core_096;
  wire cgp_core_097;

  assign cgp_core_018 = ~input_a[1];
  assign cgp_core_019 = input_a[1] & input_c[0];
  assign cgp_core_020 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_022 = cgp_core_020 ^ cgp_core_019;
  assign cgp_core_023 = cgp_core_020 & cgp_core_019;
  assign cgp_core_025 = input_a[0] ^ cgp_core_018;
  assign cgp_core_026 = ~(input_a[0] & input_h[1]);
  assign cgp_core_028 = input_a[1] & cgp_core_022;
  assign cgp_core_034 = ~(input_g[0] & input_h[0]);
  assign cgp_core_036 = ~(input_g[1] | input_h[1]);
  assign cgp_core_037 = input_e[1] & input_a[0];
  assign cgp_core_041 = input_g[0] ^ cgp_core_034;
  assign cgp_core_042 = input_d[0] & input_g[1];
  assign cgp_core_044 = input_d[0] & input_c[0];
  assign cgp_core_045_not = ~input_a[0];
  assign cgp_core_046_not = ~cgp_core_042;
  assign cgp_core_047 = ~(cgp_core_044 & input_e[1]);
  assign cgp_core_050 = ~(cgp_core_025 & input_h[1]);
  assign cgp_core_051 = cgp_core_025 & cgp_core_041;
  assign cgp_core_052_not = ~input_e[0];
  assign cgp_core_054 = input_a[1] ^ cgp_core_051;
  assign cgp_core_055 = ~cgp_core_052_not;
  assign cgp_core_056 = cgp_core_045_not | cgp_core_055;
  assign cgp_core_059 = cgp_core_047 ^ cgp_core_056;
  assign cgp_core_060 = ~cgp_core_047;
  assign cgp_core_061 = ~input_h[0];
  assign cgp_core_062 = ~(input_f[0] ^ input_a[0]);
  assign cgp_core_068 = input_e[0] & input_f[0];
  assign cgp_core_069 = input_g[1] ^ input_f[1];
  assign cgp_core_070 = input_e[1] ^ input_e[1];
  assign cgp_core_071 = input_f[1] | input_d[1];
  assign cgp_core_072 = input_c[0] & cgp_core_068;
  assign cgp_core_076 = input_f[1] | input_g[0];
  assign cgp_core_078 = input_b[1] ^ cgp_core_072;
  assign cgp_core_079 = ~(input_e[0] & cgp_core_078);
  assign cgp_core_082 = ~(input_a[1] ^ input_c[0]);
  assign cgp_core_083 = ~cgp_core_071;
  assign cgp_core_084 = ~(cgp_core_054 | input_h[1]);
  assign cgp_core_085 = ~(cgp_core_084 ^ cgp_core_082);
  assign cgp_core_088 = ~(input_e[0] | input_g[1]);
  assign cgp_core_091 = ~(cgp_core_050 ^ input_a[0]);
  assign cgp_core_094 = input_c[0] | input_a[1];
  assign cgp_core_096 = ~(input_d[1] & input_a[1]);
  assign cgp_core_097 = cgp_core_094 | cgp_core_096;

  assign cgp_out[0] = 1'b1;
endmodule