module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_066_not;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_101;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_110;

  assign cgp_core_020 = input_h[0] ^ input_a[1];
  assign cgp_core_025 = ~(input_i[0] ^ input_h[0]);
  assign cgp_core_027 = input_d[0] ^ input_h[0];
  assign cgp_core_029 = input_f[1] ^ input_e[1];
  assign cgp_core_031 = input_h[0] & input_i[1];
  assign cgp_core_032 = ~(input_g[0] ^ input_h[1]);
  assign cgp_core_033 = input_e[1] | cgp_core_032;
  assign cgp_core_034_not = ~input_e[1];
  assign cgp_core_037 = ~(input_h[0] ^ input_b[0]);
  assign cgp_core_039 = ~(input_g[1] & input_c[1]);
  assign cgp_core_040 = ~(input_c[0] ^ input_c[1]);
  assign cgp_core_042 = cgp_core_039 ^ input_c[0];
  assign cgp_core_043 = ~(input_a[0] & input_a[1]);
  assign cgp_core_046 = input_g[0] & cgp_core_040;
  assign cgp_core_047 = input_b[0] ^ input_c[0];
  assign cgp_core_049 = ~(input_g[1] ^ input_d[1]);
  assign cgp_core_050 = input_b[1] ^ cgp_core_049;
  assign cgp_core_051 = input_e[0] ^ input_d[1];
  assign cgp_core_052 = input_b[1] ^ input_g[0];
  assign cgp_core_054 = ~(input_f[1] ^ input_g[1]);
  assign cgp_core_055 = ~(input_f[1] & input_e[0]);
  assign cgp_core_056 = ~cgp_core_054;
  assign cgp_core_057 = ~(cgp_core_054 ^ input_a[0]);
  assign cgp_core_058 = cgp_core_055 | input_i[0];
  assign cgp_core_059 = input_f[0] ^ input_g[0];
  assign cgp_core_060 = ~input_e[0];
  assign cgp_core_064 = ~input_g[1];
  assign cgp_core_066_not = ~cgp_core_058;
  assign cgp_core_069 = cgp_core_043 ^ input_i[0];
  assign cgp_core_070 = input_g[1] ^ input_i[1];
  assign cgp_core_071 = cgp_core_047 & cgp_core_060;
  assign cgp_core_073 = input_h[0] & cgp_core_069;
  assign cgp_core_074 = ~(cgp_core_071 | input_d[1]);
  assign cgp_core_075 = ~input_f[0];
  assign cgp_core_076 = input_i[0] & cgp_core_066_not;
  assign cgp_core_077 = input_i[1] ^ cgp_core_074;
  assign cgp_core_078 = input_g[1] & cgp_core_074;
  assign cgp_core_079 = ~(input_h[0] & input_g[0]);
  assign cgp_core_081 = input_d[0] | input_d[0];
  assign cgp_core_082 = input_f[0] ^ cgp_core_079;
  assign cgp_core_083 = input_b[1] & cgp_core_079;
  assign cgp_core_084 = input_g[0] | cgp_core_083;
  assign cgp_core_085 = input_g[1] & input_g[1];
  assign cgp_core_086 = ~(input_f[1] ^ input_a[1]);
  assign cgp_core_090 = ~(input_i[1] & input_h[1]);
  assign cgp_core_091 = ~input_e[0];
  assign cgp_core_092 = ~input_b[0];
  assign cgp_core_093 = input_b[1] | input_b[0];
  assign cgp_core_094 = input_d[1] & input_i[1];
  assign cgp_core_095 = ~(input_d[0] & cgp_core_077);
  assign cgp_core_096 = ~(input_g[1] | input_g[0]);
  assign cgp_core_098 = ~cgp_core_031;
  assign cgp_core_099 = input_e[1] & cgp_core_096;
  assign cgp_core_100 = ~cgp_core_031;
  assign cgp_core_101 = input_i[0] & cgp_core_096;
  assign cgp_core_106 = ~(input_f[0] & cgp_core_101);
  assign cgp_core_107 = cgp_core_099 | cgp_core_094;
  assign cgp_core_110 = input_d[1] | input_a[0];

  assign cgp_out[0] = 1'b0;
endmodule