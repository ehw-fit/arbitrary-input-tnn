module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052_not;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059_not;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;

  assign cgp_core_014 = ~input_d[1];
  assign cgp_core_016 = ~(input_a[1] & input_d[0]);
  assign cgp_core_018 = input_b[0] | input_f[0];
  assign cgp_core_020 = ~(input_a[0] & input_c[0]);
  assign cgp_core_024 = input_d[1] ^ input_c[1];
  assign cgp_core_025 = input_b[0] | input_b[0];
  assign cgp_core_026 = input_c[0] & input_b[1];
  assign cgp_core_027 = ~(input_b[1] | input_f[0]);
  assign cgp_core_029 = input_c[1] ^ input_a[0];
  assign cgp_core_031 = ~(input_d[1] ^ input_b[1]);
  assign cgp_core_034 = ~(input_e[0] | input_d[0]);
  assign cgp_core_035_not = ~input_e[1];
  assign cgp_core_037 = ~(input_f[0] ^ input_c[0]);
  assign cgp_core_038 = ~input_a[0];
  assign cgp_core_039 = input_d[0] | input_a[0];
  assign cgp_core_041 = ~(input_f[1] | input_d[0]);
  assign cgp_core_043 = input_a[0] & input_d[0];
  assign cgp_core_044 = ~input_e[0];
  assign cgp_core_046 = input_b[1] | input_e[1];
  assign cgp_core_047 = ~(input_f[0] ^ input_a[1]);
  assign cgp_core_048 = ~cgp_core_046;
  assign cgp_core_050 = input_a[1] & input_c[1];
  assign cgp_core_051 = cgp_core_050 & cgp_core_048;
  assign cgp_core_052_not = ~input_e[0];
  assign cgp_core_053 = ~(input_e[0] ^ input_b[0]);
  assign cgp_core_054 = ~input_d[0];
  assign cgp_core_056 = input_b[1] | input_c[0];
  assign cgp_core_057 = ~(input_c[0] ^ input_a[1]);
  assign cgp_core_058 = input_a[0] | input_c[0];
  assign cgp_core_059_not = ~input_e[1];
  assign cgp_core_060 = input_e[1] & input_f[1];
  assign cgp_core_061 = input_c[1] | input_a[0];
  assign cgp_core_062 = input_b[0] & input_a[0];
  assign cgp_core_065 = ~(input_a[1] ^ input_e[1]);
  assign cgp_core_066 = ~(input_d[0] ^ input_c[1]);

  assign cgp_out[0] = cgp_core_051;
endmodule