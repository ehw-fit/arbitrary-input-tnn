module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;

  assign cgp_core_017 = input_b[0] ^ input_c[0];
  assign cgp_core_018 = ~(input_b[0] | input_c[0]);
  assign cgp_core_019 = input_b[1] ^ input_e[1];
  assign cgp_core_020 = ~(input_b[1] | input_c[1]);
  assign cgp_core_021 = cgp_core_019 | input_b[0];
  assign cgp_core_022 = cgp_core_019 & input_d[2];
  assign cgp_core_023 = input_d[0] | cgp_core_022;
  assign cgp_core_024 = ~(input_b[2] | input_b[2]);
  assign cgp_core_025 = input_b[2] & input_d[1];
  assign cgp_core_026_not = ~input_c[0];
  assign cgp_core_027 = cgp_core_024 & cgp_core_023;
  assign cgp_core_028 = cgp_core_025 | input_d[0];
  assign cgp_core_029 = ~input_d[0];
  assign cgp_core_030 = input_d[0] & input_e[0];
  assign cgp_core_031 = input_b[1] ^ input_e[1];
  assign cgp_core_032 = input_c[1] & input_e[1];
  assign cgp_core_033 = input_e[1] ^ cgp_core_030;
  assign cgp_core_036 = input_d[2] & input_e[0];
  assign cgp_core_037 = ~input_d[2];
  assign cgp_core_038 = cgp_core_036 ^ input_e[0];
  assign cgp_core_039 = cgp_core_036 & input_c[0];
  assign cgp_core_043 = input_d[1] ^ cgp_core_033;
  assign cgp_core_045 = ~(cgp_core_043 & input_d[1]);
  assign cgp_core_049 = cgp_core_026_not & cgp_core_038;
  assign cgp_core_052 = ~(input_e[2] & cgp_core_026_not);
  assign cgp_core_054 = cgp_core_028 & input_e[0];
  assign cgp_core_055 = input_d[2] ^ input_b[2];
  assign cgp_core_056 = input_d[2] & cgp_core_052;
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058 = cgp_core_057 & input_e[0];
  assign cgp_core_059 = ~input_e[1];
  assign cgp_core_060 = ~cgp_core_055;
  assign cgp_core_061 = ~input_e[1];
  assign cgp_core_062 = ~(cgp_core_061 & cgp_core_059);
  assign cgp_core_063 = ~input_b[2];
  assign cgp_core_064 = input_a[2] & cgp_core_063;
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066 = ~(input_a[2] ^ input_a[0]);
  assign cgp_core_067 = input_a[0] & input_a[1];
  assign cgp_core_068 = ~input_b[0];
  assign cgp_core_069 = input_a[1] & cgp_core_068;
  assign cgp_core_070 = input_d[2] & cgp_core_067;
  assign cgp_core_071 = input_a[1] & input_e[2];
  assign cgp_core_073 = ~cgp_core_017;
  assign cgp_core_074 = input_b[0] & input_b[1];
  assign cgp_core_075 = input_c[2] & cgp_core_067;
  assign cgp_core_076 = ~(input_a[0] & input_a[0]);
  assign cgp_core_077 = cgp_core_076 & cgp_core_067;

  assign cgp_out[0] = 1'b0;
endmodule