module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;

  assign cgp_core_011 = input_a[0] ^ input_b[0];
  assign cgp_core_012 = input_a[0] & input_b[0];
  assign cgp_core_013 = input_a[1] ^ input_b[1];
  assign cgp_core_014 = ~(input_a[1] & input_b[1]);
  assign cgp_core_015 = cgp_core_013 ^ cgp_core_012;
  assign cgp_core_018 = ~(input_a[2] & input_b[2]);
  assign cgp_core_019 = input_a[2] & input_b[2];
  assign cgp_core_021 = cgp_core_018 & input_b[2];
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_023 = ~cgp_core_022;
  assign cgp_core_024 = ~input_c[2];
  assign cgp_core_025 = cgp_core_018 & cgp_core_024;
  assign cgp_core_026 = input_a[1] & cgp_core_023;
  assign cgp_core_027 = cgp_core_018 & input_c[2];
  assign cgp_core_028 = cgp_core_027 & cgp_core_023;
  assign cgp_core_029 = ~input_c[1];
  assign cgp_core_030 = cgp_core_015 & cgp_core_029;
  assign cgp_core_031 = cgp_core_030 & cgp_core_028;
  assign cgp_core_032 = ~(input_c[1] ^ input_c[1]);
  assign cgp_core_033 = cgp_core_032 & cgp_core_028;
  assign cgp_core_034 = ~input_c[0];
  assign cgp_core_035 = input_a[1] & cgp_core_034;
  assign cgp_core_036 = cgp_core_035 & cgp_core_033;
  assign cgp_core_037 = ~(cgp_core_011 ^ input_c[0]);
  assign cgp_core_038 = cgp_core_037 & cgp_core_033;
  assign cgp_core_039 = cgp_core_036 | cgp_core_031;
  assign cgp_core_040 = cgp_core_022 | input_a[0];

  assign cgp_out[0] = 1'b1;
endmodule