module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058_not;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080_not;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_091;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_021 = input_d[2] ^ input_c[1];
  assign cgp_core_022 = ~(input_d[1] ^ input_c[0]);
  assign cgp_core_023 = input_d[0] ^ input_b[1];
  assign cgp_core_025 = ~input_d[0];
  assign cgp_core_027 = input_c[2] | input_e[2];
  assign cgp_core_028 = input_c[2] & input_e[2];
  assign cgp_core_029 = input_e[1] | input_c[1];
  assign cgp_core_030 = cgp_core_027 & input_a[1];
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = input_a[2] & input_b[2];
  assign cgp_core_035 = input_f[1] & input_f[2];
  assign cgp_core_036 = input_b[2] ^ input_f[0];
  assign cgp_core_037 = ~(input_d[0] & input_e[2]);
  assign cgp_core_040 = input_a[2] & cgp_core_029;
  assign cgp_core_041 = input_a[0] | input_a[1];
  assign cgp_core_044 = cgp_core_031 | cgp_core_040;
  assign cgp_core_045 = ~(input_a[2] ^ input_b[1]);
  assign cgp_core_047 = ~(input_b[0] ^ input_c[1]);
  assign cgp_core_051 = input_a[2] | input_a[1];
  assign cgp_core_052 = ~(input_d[1] & input_d[0]);
  assign cgp_core_053 = input_f[0] | input_e[2];
  assign cgp_core_054 = input_d[2] & input_f[2];
  assign cgp_core_056 = ~(input_d[1] | input_f[0]);
  assign cgp_core_058_not = ~input_b[0];
  assign cgp_core_059 = input_a[2] ^ input_a[2];
  assign cgp_core_062 = ~(input_f[1] ^ input_c[1]);
  assign cgp_core_063 = ~(input_d[2] | input_d[2]);
  assign cgp_core_065 = ~(input_b[0] | input_f[2]);
  assign cgp_core_069 = input_c[1] & input_b[2];
  assign cgp_core_071 = cgp_core_054 & input_b[2];
  assign cgp_core_072 = input_d[1] ^ input_f[2];
  assign cgp_core_073 = input_b[2] ^ input_f[2];
  assign cgp_core_074_not = ~cgp_core_071;
  assign cgp_core_075 = ~(input_e[1] | input_f[0]);
  assign cgp_core_077 = cgp_core_044 & cgp_core_074_not;
  assign cgp_core_078 = ~(input_a[0] ^ input_b[0]);
  assign cgp_core_080_not = ~input_d[2];
  assign cgp_core_081 = ~input_d[1];
  assign cgp_core_082 = ~(input_f[2] | input_a[0]);
  assign cgp_core_083 = input_d[2] ^ input_a[0];
  assign cgp_core_086 = ~(input_d[2] & input_e[0]);
  assign cgp_core_088 = input_f[0] | input_c[1];
  assign cgp_core_089 = ~(input_b[1] | input_c[1]);
  assign cgp_core_091 = ~(input_e[2] | input_a[1]);
  assign cgp_core_094 = input_d[1] | input_f[0];
  assign cgp_core_095 = ~(input_f[0] & input_a[2]);
  assign cgp_core_098 = input_b[0] ^ input_a[2];
  assign cgp_core_099 = ~input_f[1];

  assign cgp_out[0] = cgp_core_077;
endmodule