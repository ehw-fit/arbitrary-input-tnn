module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044_not;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;

  assign cgp_core_012 = ~(input_d[1] & input_b[1]);
  assign cgp_core_014 = ~(input_e[0] ^ input_e[0]);
  assign cgp_core_015 = input_a[0] ^ input_a[1];
  assign cgp_core_016 = ~input_b[1];
  assign cgp_core_018 = input_e[1] | input_b[1];
  assign cgp_core_022 = input_d[1] & input_a[1];
  assign cgp_core_023 = input_c[0] & input_b[1];
  assign cgp_core_024 = ~(input_a[0] | input_a[1]);
  assign cgp_core_025 = ~(input_d[1] & input_d[1]);
  assign cgp_core_026 = cgp_core_018 | input_a[1];
  assign cgp_core_027 = input_e[1] & input_a[1];
  assign cgp_core_030 = ~(input_d[0] | input_b[0]);
  assign cgp_core_031 = input_c[1] & input_d[1];
  assign cgp_core_032 = ~input_d[1];
  assign cgp_core_033 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_035 = ~input_b[1];
  assign cgp_core_036 = ~cgp_core_031;
  assign cgp_core_037 = cgp_core_026 & cgp_core_036;
  assign cgp_core_041 = ~(input_c[0] ^ input_e[1]);
  assign cgp_core_042 = ~(input_e[1] & input_e[0]);
  assign cgp_core_043 = ~(input_b[1] & input_c[1]);
  assign cgp_core_044_not = ~input_e[0];
  assign cgp_core_045 = ~(input_b[0] & input_c[1]);
  assign cgp_core_046 = input_b[1] & input_e[1];
  assign cgp_core_047 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_048 = input_b[1] | input_a[1];
  assign cgp_core_049 = input_a[1] | input_b[0];
  assign cgp_core_051 = ~(input_d[1] ^ input_d[0]);
  assign cgp_core_053 = cgp_core_037 | cgp_core_027;

  assign cgp_out[0] = cgp_core_053;
endmodule