module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063_not;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;

  assign cgp_core_016 = ~(input_a[9] & input_a[2]);
  assign cgp_core_021 = ~(input_a[3] & input_a[0]);
  assign cgp_core_023 = input_a[5] & input_a[8];
  assign cgp_core_024 = ~(input_a[2] | input_a[6]);
  assign cgp_core_025_not = ~input_a[1];
  assign cgp_core_027 = input_a[1] | input_a[8];
  assign cgp_core_028 = input_a[12] ^ input_a[5];
  assign cgp_core_029 = ~input_a[7];
  assign cgp_core_031 = ~(input_a[12] | input_a[9]);
  assign cgp_core_033 = ~(input_a[9] ^ input_a[4]);
  assign cgp_core_034_not = ~input_a[13];
  assign cgp_core_035 = ~(input_a[13] & input_a[7]);
  assign cgp_core_037 = input_a[3] & input_a[13];
  assign cgp_core_038 = ~(input_a[3] | input_a[13]);
  assign cgp_core_040 = ~(input_a[4] ^ input_a[10]);
  assign cgp_core_045 = ~(input_a[13] | input_a[13]);
  assign cgp_core_046 = ~(input_a[10] ^ input_a[11]);
  assign cgp_core_047 = ~input_a[8];
  assign cgp_core_050 = ~(input_a[10] ^ input_a[9]);
  assign cgp_core_051 = ~input_a[3];
  assign cgp_core_055 = ~input_a[1];
  assign cgp_core_056 = input_a[10] ^ input_a[6];
  assign cgp_core_059 = input_a[3] | input_a[10];
  assign cgp_core_060 = ~input_a[2];
  assign cgp_core_061 = ~input_a[3];
  assign cgp_core_063_not = ~input_a[12];
  assign cgp_core_064 = input_a[11] & input_a[1];
  assign cgp_core_067 = ~(input_a[2] ^ input_a[3]);
  assign cgp_core_072 = input_a[0] & input_a[9];
  assign cgp_core_074 = input_a[11] | input_a[3];
  assign cgp_core_076 = ~(input_a[12] & input_a[0]);
  assign cgp_core_077 = input_a[6] ^ input_a[9];
  assign cgp_core_079 = input_a[1] | input_a[6];
  assign cgp_core_081 = ~(input_a[2] & input_a[4]);
  assign cgp_core_083 = input_a[3] & input_a[3];
  assign cgp_core_086 = input_a[7] & input_a[10];
  assign cgp_core_087 = input_a[12] & input_a[0];
  assign cgp_core_089 = input_a[5] | input_a[3];
  assign cgp_core_090 = ~(input_a[11] & input_a[0]);

  assign cgp_out[0] = 1'b0;
  assign cgp_out[1] = input_a[2];
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = 1'b0;
endmodule