module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_059_not;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_089;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_097;
  wire cgp_core_099;

  assign cgp_core_020 = input_f[0] ^ input_a[2];
  assign cgp_core_023 = input_b[2] | input_e[0];
  assign cgp_core_024 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_026 = ~(input_c[2] | input_f[2]);
  assign cgp_core_028 = ~(input_d[0] | input_a[0]);
  assign cgp_core_032_not = ~input_d[2];
  assign cgp_core_033 = ~(input_a[0] | input_c[0]);
  assign cgp_core_035 = ~input_f[1];
  assign cgp_core_037 = input_d[0] | input_b[1];
  assign cgp_core_038 = input_c[1] ^ input_e[1];
  assign cgp_core_039 = ~input_e[0];
  assign cgp_core_040 = ~input_a[1];
  assign cgp_core_042 = ~(input_b[0] & input_b[2]);
  assign cgp_core_044 = input_e[1] | input_b[2];
  assign cgp_core_046 = input_d[0] ^ input_e[1];
  assign cgp_core_048 = input_c[2] & input_d[2];
  assign cgp_core_049 = ~(input_c[0] ^ input_a[2]);
  assign cgp_core_051 = input_b[1] & input_d[2];
  assign cgp_core_052 = input_a[1] | input_d[0];
  assign cgp_core_053 = ~input_a[2];
  assign cgp_core_055 = ~input_d[2];
  assign cgp_core_057 = ~(input_f[2] ^ input_b[2]);
  assign cgp_core_059_not = ~input_d[2];
  assign cgp_core_061 = ~(input_c[2] | input_a[2]);
  assign cgp_core_062 = ~(input_f[0] ^ input_f[0]);
  assign cgp_core_063 = ~input_e[1];
  assign cgp_core_065 = ~input_f[1];
  assign cgp_core_066 = ~(input_b[1] ^ input_e[2]);
  assign cgp_core_068 = ~input_f[0];
  assign cgp_core_069_not = ~input_f[2];
  assign cgp_core_072 = input_d[0] & input_a[0];
  assign cgp_core_075 = ~input_d[2];
  assign cgp_core_076 = input_a[2] & cgp_core_075;
  assign cgp_core_078 = ~(input_c[2] | input_d[0]);
  assign cgp_core_079 = ~(input_d[0] & input_a[2]);
  assign cgp_core_082 = input_a[0] & input_c[1];
  assign cgp_core_083 = ~(input_e[0] ^ input_b[0]);
  assign cgp_core_089 = input_a[1] ^ input_c[0];
  assign cgp_core_092 = input_e[2] & input_c[2];
  assign cgp_core_093 = ~input_a[1];
  assign cgp_core_094 = ~input_a[1];
  assign cgp_core_097 = ~(input_f[0] ^ input_b[1]);
  assign cgp_core_099 = cgp_core_092 | cgp_core_076;

  assign cgp_out[0] = cgp_core_099;
endmodule