module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075_not;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_094;
  wire cgp_core_095;

  assign cgp_core_019 = input_b[0] ^ input_c[0];
  assign cgp_core_020 = input_b[1] ^ input_c[0];
  assign cgp_core_021 = input_d[0] & input_e[1];
  assign cgp_core_022 = ~(input_g[0] | cgp_core_019);
  assign cgp_core_023 = cgp_core_020 & cgp_core_019;
  assign cgp_core_024 = cgp_core_021 | input_f[1];
  assign cgp_core_025 = input_d[0] ^ input_c[0];
  assign cgp_core_026 = ~(input_a[0] & input_h[0]);
  assign cgp_core_027 = ~(input_a[1] | input_a[1]);
  assign cgp_core_028 = input_a[1] & input_d[1];
  assign cgp_core_029 = cgp_core_027 ^ cgp_core_026;
  assign cgp_core_030 = input_b[1] & input_f[1];
  assign cgp_core_031 = input_c[1] | cgp_core_030;
  assign cgp_core_032 = input_c[0] ^ cgp_core_031;
  assign cgp_core_033 = input_a[1] & input_f[1];
  assign cgp_core_034 = input_g[0] ^ input_h[0];
  assign cgp_core_035 = input_g[0] & input_h[0];
  assign cgp_core_036 = input_g[1] & input_h[1];
  assign cgp_core_037 = input_g[1] & input_h[1];
  assign cgp_core_038 = ~cgp_core_036;
  assign cgp_core_039 = cgp_core_036 & cgp_core_035;
  assign cgp_core_040 = input_f[1] | input_b[1];
  assign cgp_core_041 = input_e[1] ^ input_b[1];
  assign cgp_core_042 = input_d[0] & input_e[0];
  assign cgp_core_043 = input_d[1] & cgp_core_038;
  assign cgp_core_044 = input_b[1] & cgp_core_038;
  assign cgp_core_046 = cgp_core_043 & input_f[1];
  assign cgp_core_047 = ~(cgp_core_044 | cgp_core_046);
  assign cgp_core_048 = input_a[0] ^ cgp_core_047;
  assign cgp_core_049 = ~cgp_core_040;
  assign cgp_core_050 = ~(input_c[0] & input_d[1]);
  assign cgp_core_051 = ~(cgp_core_025 | cgp_core_041);
  assign cgp_core_052 = ~(input_e[1] & input_f[0]);
  assign cgp_core_053 = cgp_core_029 & input_f[0];
  assign cgp_core_054 = cgp_core_052 | cgp_core_051;
  assign cgp_core_056 = input_c[0] | input_c[1];
  assign cgp_core_057 = ~(cgp_core_032 | cgp_core_048);
  assign cgp_core_058 = cgp_core_032 & cgp_core_048;
  assign cgp_core_059 = input_a[1] ^ cgp_core_056;
  assign cgp_core_060 = cgp_core_057 & cgp_core_056;
  assign cgp_core_061 = ~(cgp_core_058 | cgp_core_060);
  assign cgp_core_063 = cgp_core_033 & cgp_core_049;
  assign cgp_core_064_not = ~cgp_core_061;
  assign cgp_core_067 = input_e[0] ^ input_f[0];
  assign cgp_core_068 = input_e[0] & input_d[0];
  assign cgp_core_069 = input_c[0] ^ input_f[1];
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = input_a[0] | cgp_core_072;
  assign cgp_core_074 = ~(input_a[1] | input_a[1]);
  assign cgp_core_075_not = ~cgp_core_074;
  assign cgp_core_076 = ~cgp_core_064_not;
  assign cgp_core_077 = input_g[1] & input_a[0];
  assign cgp_core_078 = input_c[0] ^ input_c[1];
  assign cgp_core_079 = input_f[0] & cgp_core_078;
  assign cgp_core_080 = cgp_core_079 & input_h[0];
  assign cgp_core_081 = ~(cgp_core_059 ^ cgp_core_073);
  assign cgp_core_082 = cgp_core_081 & input_b[1];
  assign cgp_core_083 = ~cgp_core_071;
  assign cgp_core_084 = input_g[0] & cgp_core_083;
  assign cgp_core_089 = input_a[0] & cgp_core_067;
  assign cgp_core_090 = input_a[0] & input_c[0];
  assign cgp_core_091 = ~(cgp_core_050 ^ input_f[1]);
  assign cgp_core_094 = ~(cgp_core_090 & input_c[0]);
  assign cgp_core_095 = ~input_a[1];

  assign cgp_out[0] = 1'b1;
endmodule