module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_021_not;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_075;
  wire cgp_core_076_not;
  wire cgp_core_078;
  wire cgp_core_079_not;
  wire cgp_core_080_not;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_090;

  assign cgp_core_018 = ~(input_a[8] | input_a[9]);
  assign cgp_core_021_not = ~input_a[2];
  assign cgp_core_022 = ~(input_a[7] & input_a[2]);
  assign cgp_core_023 = ~(input_a[10] | input_a[8]);
  assign cgp_core_025 = input_a[1] | input_a[7];
  assign cgp_core_026 = input_a[11] | input_a[11];
  assign cgp_core_027 = input_a[9] ^ input_a[1];
  assign cgp_core_029 = input_a[9] & input_a[0];
  assign cgp_core_033 = ~input_a[13];
  assign cgp_core_034 = ~(input_a[13] ^ input_a[10]);
  assign cgp_core_035 = input_a[12] | input_a[3];
  assign cgp_core_037 = ~input_a[10];
  assign cgp_core_041 = input_a[1] ^ input_a[0];
  assign cgp_core_042 = input_a[10] & input_a[8];
  assign cgp_core_048 = ~(input_a[7] & input_a[2]);
  assign cgp_core_050 = ~(input_a[8] | input_a[2]);
  assign cgp_core_052 = input_a[11] | input_a[8];
  assign cgp_core_053 = ~(input_a[12] & input_a[4]);
  assign cgp_core_054 = ~input_a[9];
  assign cgp_core_056 = input_a[0] & input_a[10];
  assign cgp_core_059 = input_a[1] & input_a[9];
  assign cgp_core_060 = ~(input_a[3] ^ input_a[5]);
  assign cgp_core_064 = ~(input_a[12] ^ input_a[5]);
  assign cgp_core_065 = ~(input_a[2] | input_a[7]);
  assign cgp_core_067 = input_a[13] | input_a[5];
  assign cgp_core_070 = input_a[12] ^ input_a[3];
  assign cgp_core_071 = ~input_a[6];
  assign cgp_core_075 = input_a[3] | input_a[0];
  assign cgp_core_076_not = ~input_a[9];
  assign cgp_core_078 = ~(input_a[3] ^ input_a[0]);
  assign cgp_core_079_not = ~input_a[12];
  assign cgp_core_080_not = ~input_a[12];
  assign cgp_core_081 = ~input_a[12];
  assign cgp_core_082 = ~(input_a[2] ^ input_a[2]);
  assign cgp_core_084 = ~(input_a[11] | input_a[4]);
  assign cgp_core_085 = ~(input_a[9] | input_a[13]);
  assign cgp_core_086 = ~(input_a[9] ^ input_a[6]);
  assign cgp_core_088 = ~(input_a[3] ^ input_a[1]);
  assign cgp_core_090 = ~input_a[4];

  assign cgp_out[0] = input_a[13];
  assign cgp_out[1] = 1'b1;
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = 1'b0;
endmodule