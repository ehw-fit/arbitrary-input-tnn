module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039_not;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;

  assign cgp_core_012 = ~input_c[0];
  assign cgp_core_013 = input_b[0] & input_b[1];
  assign cgp_core_015 = input_c[0] & input_b[1];
  assign cgp_core_016 = input_e[1] ^ input_a[0];
  assign cgp_core_017 = ~(input_e[1] | input_b[1]);
  assign cgp_core_018 = ~input_c[0];
  assign cgp_core_019 = input_c[1] | input_c[0];
  assign cgp_core_021 = input_a[0] | input_b[1];
  assign cgp_core_024_not = ~input_d[1];
  assign cgp_core_025 = input_e[0] | input_e[1];
  assign cgp_core_026 = ~(input_e[1] & input_c[0]);
  assign cgp_core_027 = input_a[1] & cgp_core_025;
  assign cgp_core_029 = ~(input_d[0] ^ input_a[0]);
  assign cgp_core_031 = input_c[1] & input_d[1];
  assign cgp_core_033 = ~(input_d[1] ^ input_a[0]);
  assign cgp_core_035_not = ~input_a[1];
  assign cgp_core_036 = ~(input_b[0] & input_d[1]);
  assign cgp_core_037 = ~(input_b[1] | input_d[1]);
  assign cgp_core_038 = ~(input_a[1] & input_e[0]);
  assign cgp_core_039_not = ~cgp_core_031;
  assign cgp_core_041 = ~(input_b[0] & input_e[0]);
  assign cgp_core_043 = cgp_core_021 & cgp_core_039_not;
  assign cgp_core_045 = input_c[0] ^ input_b[1];
  assign cgp_core_046 = ~input_c[0];
  assign cgp_core_050 = input_e[1] & input_b[0];
  assign cgp_core_052 = cgp_core_027 | cgp_core_050;
  assign cgp_core_054 = cgp_core_043 | cgp_core_052;

  assign cgp_out[0] = cgp_core_054;
endmodule