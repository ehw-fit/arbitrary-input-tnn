module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_096;
  wire cgp_core_097;

  assign cgp_core_021 = input_g[1] | input_d[1];
  assign cgp_core_022 = ~(input_e[0] & input_b[0]);
  assign cgp_core_023 = input_e[0] & input_e[1];
  assign cgp_core_024 = ~(input_h[0] ^ cgp_core_023);
  assign cgp_core_025_not = ~input_a[0];
  assign cgp_core_026_not = ~input_c[0];
  assign cgp_core_027 = input_a[1] ^ input_d[1];
  assign cgp_core_029 = ~cgp_core_027;
  assign cgp_core_030 = ~(cgp_core_027 & input_h[0]);
  assign cgp_core_031 = input_a[0] & input_f[1];
  assign cgp_core_032 = ~(input_a[1] ^ input_c[1]);
  assign cgp_core_033 = input_e[0] & input_b[1];
  assign cgp_core_034 = ~(input_g[0] & input_b[0]);
  assign cgp_core_035 = input_e[1] & input_g[1];
  assign cgp_core_037 = input_b[0] & input_h[1];
  assign cgp_core_039 = input_e[1] ^ cgp_core_035;
  assign cgp_core_040 = cgp_core_037 | input_h[1];
  assign cgp_core_043 = input_g[0] ^ input_c[1];
  assign cgp_core_045 = input_d[1] & input_c[0];
  assign cgp_core_046 = ~(cgp_core_043 ^ input_g[1]);
  assign cgp_core_050 = input_e[1] ^ input_f[1];
  assign cgp_core_051 = ~(input_d[1] | input_g[0]);
  assign cgp_core_053 = cgp_core_029 & input_g[1];
  assign cgp_core_054 = ~(input_g[1] & cgp_core_051);
  assign cgp_core_055 = ~(input_b[1] & cgp_core_051);
  assign cgp_core_056 = input_d[0] | input_g[1];
  assign cgp_core_058 = input_g[1] | input_a[1];
  assign cgp_core_060 = ~(input_c[0] ^ input_b[1]);
  assign cgp_core_061 = ~(input_h[1] & input_a[1]);
  assign cgp_core_062 = input_h[0] ^ input_c[1];
  assign cgp_core_064_not = ~cgp_core_061;
  assign cgp_core_065 = ~input_e[1];
  assign cgp_core_067 = ~(input_e[0] & input_h[0]);
  assign cgp_core_069 = input_a[0] | input_e[0];
  assign cgp_core_070 = ~(input_e[1] | input_c[1]);
  assign cgp_core_072 = input_a[1] ^ input_g[1];
  assign cgp_core_073 = ~input_c[1];
  assign cgp_core_076 = ~(cgp_core_064_not | input_d[0]);
  assign cgp_core_077 = cgp_core_076 & input_d[0];
  assign cgp_core_078 = ~input_g[1];
  assign cgp_core_080 = ~(input_e[0] ^ cgp_core_077);
  assign cgp_core_082 = ~(input_g[0] ^ input_f[1]);
  assign cgp_core_084 = input_g[1] ^ input_d[0];
  assign cgp_core_085 = input_f[0] | input_b[1];
  assign cgp_core_086 = input_b[0] ^ input_a[0];
  assign cgp_core_091 = ~(cgp_core_050 ^ input_g[0]);
  assign cgp_core_092 = input_d[0] & input_a[0];
  assign cgp_core_096 = ~input_a[1];
  assign cgp_core_097 = input_c[1] | input_h[0];

  assign cgp_out[0] = 1'b1;
endmodule