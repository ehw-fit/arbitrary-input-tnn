module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_039_not;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_052;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_076;

  assign cgp_core_018 = ~(input_b[0] & input_e[1]);
  assign cgp_core_019 = input_c[2] ^ input_e[1];
  assign cgp_core_020 = input_d[2] ^ input_c[1];
  assign cgp_core_021 = ~input_d[0];
  assign cgp_core_025 = ~(input_b[0] | input_a[1]);
  assign cgp_core_026 = ~input_c[1];
  assign cgp_core_028 = cgp_core_025 | input_e[2];
  assign cgp_core_030 = ~(input_d[0] & input_b[2]);
  assign cgp_core_031 = ~(input_d[1] | input_b[0]);
  assign cgp_core_033 = cgp_core_031 ^ cgp_core_030;
  assign cgp_core_034 = input_e[2] & input_a[1];
  assign cgp_core_036 = ~(input_c[1] & input_e[2]);
  assign cgp_core_037 = input_b[0] & input_c[1];
  assign cgp_core_039_not = ~cgp_core_036;
  assign cgp_core_040 = input_c[2] | input_e[0];
  assign cgp_core_044 = ~(input_c[0] | input_e[1]);
  assign cgp_core_045 = input_a[0] ^ input_c[2];
  assign cgp_core_047 = ~(input_b[1] ^ input_e[2]);
  assign cgp_core_049 = input_e[1] | input_d[2];
  assign cgp_core_050_not = ~cgp_core_047;
  assign cgp_core_052 = cgp_core_049 | input_e[0];
  assign cgp_core_053_not = ~cgp_core_040;
  assign cgp_core_054 = cgp_core_028 & cgp_core_040;
  assign cgp_core_055 = ~(cgp_core_053_not ^ input_b[2]);
  assign cgp_core_059 = ~cgp_core_054;
  assign cgp_core_060 = ~cgp_core_055;
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_063 = input_e[0] & cgp_core_050_not;
  assign cgp_core_064 = input_d[2] | input_c[1];
  assign cgp_core_066 = ~(input_a[1] ^ input_c[1]);
  assign cgp_core_068 = ~input_a[2];
  assign cgp_core_069 = input_a[1] & input_a[2];
  assign cgp_core_070 = cgp_core_069 & input_c[2];
  assign cgp_core_071 = input_a[1] ^ input_d[1];
  assign cgp_core_076 = ~input_a[0];

  assign cgp_out[0] = 1'b0;
endmodule