module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_014_not;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_038_not;
  wire cgp_core_039_not;
  wire cgp_core_042;

  assign cgp_core_012 = input_b[2] | input_a[1];
  assign cgp_core_014_not = ~input_a[0];
  assign cgp_core_015 = input_b[1] & input_b[1];
  assign cgp_core_016 = input_a[1] ^ input_a[1];
  assign cgp_core_018 = input_a[2] | input_c[2];
  assign cgp_core_019 = input_a[2] & input_c[2];
  assign cgp_core_021 = ~(input_a[1] ^ input_a[2]);
  assign cgp_core_022 = cgp_core_019 | input_c[1];
  assign cgp_core_023 = ~(input_c[0] | input_a[0]);
  assign cgp_core_024 = ~cgp_core_022;
  assign cgp_core_025 = ~cgp_core_018;
  assign cgp_core_026 = input_b[2] & cgp_core_025;
  assign cgp_core_028 = ~input_a[0];
  assign cgp_core_029 = input_b[2] & cgp_core_024;
  assign cgp_core_032 = input_b[1] & cgp_core_029;
  assign cgp_core_036 = input_c[1] | input_b[0];
  assign cgp_core_038_not = ~input_a[0];
  assign cgp_core_039_not = ~input_a[1];
  assign cgp_core_042 = cgp_core_032 | cgp_core_026;

  assign cgp_out[0] = cgp_core_042;
endmodule