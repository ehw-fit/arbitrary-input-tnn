module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_047_not;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073_not;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_088;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_099;

  assign cgp_core_020 = ~(input_b[2] ^ input_b[2]);
  assign cgp_core_021 = ~(input_c[2] | input_d[0]);
  assign cgp_core_022 = input_f[1] & input_c[0];
  assign cgp_core_024 = input_b[1] | input_c[0];
  assign cgp_core_026 = ~(input_f[2] | input_b[0]);
  assign cgp_core_027 = input_c[0] ^ input_e[1];
  assign cgp_core_028 = input_d[1] ^ input_e[2];
  assign cgp_core_030 = input_c[2] | input_c[0];
  assign cgp_core_032 = ~input_e[2];
  assign cgp_core_036 = input_e[0] & input_f[1];
  assign cgp_core_037 = ~(input_a[0] | input_b[0]);
  assign cgp_core_038 = ~input_e[2];
  assign cgp_core_039 = ~(input_e[2] | input_c[1]);
  assign cgp_core_040 = ~input_c[1];
  assign cgp_core_043 = ~(input_e[2] ^ input_a[1]);
  assign cgp_core_045 = ~(input_b[0] ^ input_d[2]);
  assign cgp_core_047_not = ~input_a[1];
  assign cgp_core_048 = ~(input_c[1] ^ input_d[2]);
  assign cgp_core_049 = ~input_c[0];
  assign cgp_core_050 = ~(input_b[0] | input_d[0]);
  assign cgp_core_051 = ~(input_f[1] | input_c[2]);
  assign cgp_core_052 = ~input_e[1];
  assign cgp_core_053 = ~input_d[2];
  assign cgp_core_055 = input_a[1] & input_d[2];
  assign cgp_core_056 = input_d[2] & input_b[2];
  assign cgp_core_057 = input_f[2] | cgp_core_056;
  assign cgp_core_058 = ~input_a[1];
  assign cgp_core_059 = input_d[1] ^ input_a[1];
  assign cgp_core_062 = ~(input_b[0] | input_a[0]);
  assign cgp_core_065 = ~(input_c[2] ^ input_d[0]);
  assign cgp_core_066 = ~(input_d[2] | input_e[1]);
  assign cgp_core_067 = ~input_d[2];
  assign cgp_core_068 = ~(input_a[0] ^ input_c[0]);
  assign cgp_core_069 = ~input_a[1];
  assign cgp_core_070 = ~input_a[1];
  assign cgp_core_072 = ~cgp_core_057;
  assign cgp_core_073_not = ~input_d[1];
  assign cgp_core_076 = ~(input_c[0] & input_f[0]);
  assign cgp_core_077 = input_b[1] ^ input_e[0];
  assign cgp_core_079 = ~(input_f[2] ^ input_f[1]);
  assign cgp_core_081 = ~input_b[0];
  assign cgp_core_083 = ~(input_d[0] & input_a[2]);
  assign cgp_core_084 = ~(input_c[2] & input_f[0]);
  assign cgp_core_088 = input_c[0] ^ input_d[0];
  assign cgp_core_091 = ~(input_f[0] ^ input_d[2]);
  assign cgp_core_092 = input_c[0] | input_e[1];
  assign cgp_core_093 = ~input_b[2];
  assign cgp_core_096 = ~(input_c[0] | input_a[0]);
  assign cgp_core_097 = input_b[0] | input_b[0];
  assign cgp_core_099 = input_f[2] & input_f[1];

  assign cgp_out[0] = cgp_core_072;
endmodule