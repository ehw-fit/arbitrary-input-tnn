module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037_not;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063_not;
  wire cgp_core_068;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_078_not;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;

  assign cgp_core_020 = ~(input_a[0] & input_a[2]);
  assign cgp_core_022 = input_c[0] ^ input_b[1];
  assign cgp_core_023 = ~(input_a[1] | input_b[1]);
  assign cgp_core_024 = ~(input_f[0] | input_a[0]);
  assign cgp_core_025 = input_c[2] ^ input_a[0];
  assign cgp_core_026 = cgp_core_023 ^ cgp_core_025;
  assign cgp_core_027 = input_a[2] ^ input_b[1];
  assign cgp_core_028_not = ~input_a[2];
  assign cgp_core_029 = cgp_core_027 ^ input_b[2];
  assign cgp_core_032 = input_c[0] ^ input_b[1];
  assign cgp_core_033 = ~(input_f[1] ^ input_d[0]);
  assign cgp_core_034 = input_c[1] & input_b[2];
  assign cgp_core_037_not = ~cgp_core_033;
  assign cgp_core_040 = input_d[1] & input_d[0];
  assign cgp_core_044 = ~(input_f[2] | input_f[0]);
  assign cgp_core_046 = ~(input_e[1] & input_a[1]);
  assign cgp_core_047 = ~(input_b[2] & input_f[1]);
  assign cgp_core_048 = input_f[1] ^ input_e[2];
  assign cgp_core_051 = input_a[2] ^ input_f[2];
  assign cgp_core_052 = ~(input_e[2] | input_f[2]);
  assign cgp_core_054 = ~(cgp_core_051 | input_a[2]);
  assign cgp_core_055 = ~(input_c[0] & input_c[0]);
  assign cgp_core_056 = cgp_core_032 ^ cgp_core_044;
  assign cgp_core_058 = cgp_core_033 ^ cgp_core_048;
  assign cgp_core_059 = ~(input_f[2] | cgp_core_048);
  assign cgp_core_061 = input_a[2] & input_c[0];
  assign cgp_core_062 = ~(cgp_core_059 | cgp_core_061);
  assign cgp_core_063_not = ~input_a[2];
  assign cgp_core_068 = input_c[2] ^ input_b[0];
  assign cgp_core_071 = input_c[1] & input_d[1];
  assign cgp_core_072 = ~input_f[0];
  assign cgp_core_073 = ~cgp_core_072;
  assign cgp_core_074 = ~input_e[1];
  assign cgp_core_078_not = ~input_f[1];
  assign cgp_core_079 = cgp_core_078_not ^ input_d[2];
  assign cgp_core_080 = ~input_f[1];
  assign cgp_core_081 = ~(input_f[1] | cgp_core_080);
  assign cgp_core_087 = input_a[1] & input_b[0];
  assign cgp_core_088 = ~input_f[0];
  assign cgp_core_089 = cgp_core_088 & cgp_core_079;
  assign cgp_core_090 = cgp_core_056 ^ cgp_core_056;
  assign cgp_core_091 = cgp_core_020 & input_d[1];
  assign cgp_core_092 = ~cgp_core_091;
  assign cgp_core_093 = ~(cgp_core_020 ^ input_e[2]);
  assign cgp_core_094 = ~input_d[0];
  assign cgp_core_095 = input_f[1] | input_d[0];
  assign cgp_core_096 = input_b[2] | cgp_core_095;
  assign cgp_core_097 = input_d[1] | input_f[1];
  assign cgp_core_098 = ~(cgp_core_096 & cgp_core_097);

  assign cgp_out[0] = input_a[2];
endmodule