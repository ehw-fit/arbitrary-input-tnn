module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_034_not;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058_not;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067_not;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;

  assign cgp_core_017 = input_c[0] ^ input_e[0];
  assign cgp_core_020 = input_c[1] & input_e[1];
  assign cgp_core_024 = input_c[1] & input_c[0];
  assign cgp_core_025 = input_a[2] & input_e[2];
  assign cgp_core_026_not = ~input_b[1];
  assign cgp_core_029 = input_b[0] ^ cgp_core_017;
  assign cgp_core_030 = input_b[0] | cgp_core_017;
  assign cgp_core_034_not = ~input_b[0];
  assign cgp_core_037 = input_b[2] & cgp_core_026_not;
  assign cgp_core_038 = cgp_core_026_not | input_c[2];
  assign cgp_core_039 = cgp_core_026_not & input_c[2];
  assign cgp_core_040 = cgp_core_037 ^ cgp_core_039;
  assign cgp_core_041 = cgp_core_025 ^ cgp_core_040;
  assign cgp_core_042 = cgp_core_025 ^ cgp_core_040;
  assign cgp_core_043 = input_a[0] ^ input_d[0];
  assign cgp_core_044 = input_d[0] & input_d[1];
  assign cgp_core_045 = input_b[1] ^ input_d[1];
  assign cgp_core_046 = input_a[1] & input_b[1];
  assign cgp_core_047 = cgp_core_045 ^ cgp_core_044;
  assign cgp_core_048 = input_b[0] & cgp_core_044;
  assign cgp_core_049 = input_e[2] | input_d[0];
  assign cgp_core_050 = input_a[2] ^ input_d[2];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_052 = ~cgp_core_050;
  assign cgp_core_053 = cgp_core_050 & cgp_core_049;
  assign cgp_core_054 = cgp_core_051 | input_b[0];
  assign cgp_core_055 = ~cgp_core_042;
  assign cgp_core_056 = ~(cgp_core_054 & cgp_core_054);
  assign cgp_core_057 = cgp_core_041 & input_b[1];
  assign cgp_core_058_not = ~cgp_core_057;
  assign cgp_core_059 = ~(cgp_core_041 ^ input_a[2]);
  assign cgp_core_060 = ~(input_b[1] ^ cgp_core_055);
  assign cgp_core_061 = ~cgp_core_052;
  assign cgp_core_064 = ~(input_d[2] & cgp_core_052);
  assign cgp_core_065 = cgp_core_064 & cgp_core_060;
  assign cgp_core_066 = ~cgp_core_047;
  assign cgp_core_067_not = ~input_e[2];
  assign cgp_core_068 = cgp_core_067_not & cgp_core_065;
  assign cgp_core_070 = input_b[1] & cgp_core_065;
  assign cgp_core_071 = ~(cgp_core_043 | input_a[2]);
  assign cgp_core_072 = cgp_core_029 & input_c[0];
  assign cgp_core_073 = cgp_core_072 & cgp_core_070;
  assign cgp_core_076 = input_e[2] ^ cgp_core_060;

  assign cgp_out[0] = 1'b1;
endmodule