module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019_not;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036_not;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_083;

  assign cgp_core_016 = input_d[1] ^ input_a[0];
  assign cgp_core_017 = ~(input_c[1] ^ input_a[0]);
  assign cgp_core_019_not = ~input_b[1];
  assign cgp_core_023 = ~input_g[1];
  assign cgp_core_027 = ~input_a[0];
  assign cgp_core_028 = input_a[1] ^ input_f[0];
  assign cgp_core_029 = input_a[1] | input_a[0];
  assign cgp_core_030 = input_f[0] & input_a[0];
  assign cgp_core_032 = ~(input_g[1] | input_d[0]);
  assign cgp_core_035 = ~(input_g[1] | input_d[0]);
  assign cgp_core_036_not = ~input_a[1];
  assign cgp_core_038 = ~input_f[1];
  assign cgp_core_040 = ~(input_c[1] & input_c[0]);
  assign cgp_core_043 = input_a[0] ^ input_e[1];
  assign cgp_core_046 = input_f[0] & input_a[0];
  assign cgp_core_047_not = ~input_b[0];
  assign cgp_core_049 = input_g[1] | input_a[0];
  assign cgp_core_050 = input_e[1] | input_c[1];
  assign cgp_core_051 = input_g[1] | cgp_core_050;
  assign cgp_core_053 = ~input_a[1];
  assign cgp_core_054 = input_f[0] ^ input_f[1];
  assign cgp_core_055 = ~(input_d[0] & input_g[0]);
  assign cgp_core_056 = ~(input_a[0] ^ input_f[1]);
  assign cgp_core_057 = input_d[1] | input_b[1];
  assign cgp_core_058 = input_f[1] | input_f[1];
  assign cgp_core_060 = ~(input_b[1] ^ input_d[0]);
  assign cgp_core_064_not = ~input_a[0];
  assign cgp_core_065 = ~(input_d[0] & input_f[1]);
  assign cgp_core_066 = ~(input_e[0] & input_f[0]);
  assign cgp_core_067 = ~input_d[0];
  assign cgp_core_068 = ~(input_f[0] & input_e[1]);
  assign cgp_core_069 = ~(input_d[1] | input_c[1]);
  assign cgp_core_074 = ~input_c[1];
  assign cgp_core_075 = input_a[0] ^ input_f[0];
  assign cgp_core_077 = input_f[1] & input_c[1];
  assign cgp_core_078 = ~input_d[0];
  assign cgp_core_079 = ~(input_c[1] & input_d[1]);
  assign cgp_core_080 = input_d[1] | input_a[1];
  assign cgp_core_081 = input_g[0] ^ input_b[1];
  assign cgp_core_083 = cgp_core_080 | cgp_core_051;

  assign cgp_out[0] = cgp_core_083;
endmodule