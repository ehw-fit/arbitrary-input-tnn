module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048_not;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053_not;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_020 = input_f[1] ^ input_e[0];
  assign cgp_core_024 = input_d[0] ^ input_b[1];
  assign cgp_core_025 = input_a[2] & input_e[1];
  assign cgp_core_026 = ~(input_a[2] & input_b[2]);
  assign cgp_core_029 = input_b[2] & input_c[2];
  assign cgp_core_030 = input_b[0] & input_f[0];
  assign cgp_core_031 = input_b[0] & input_b[0];
  assign cgp_core_033 = ~(input_d[2] & input_a[0]);
  assign cgp_core_034 = input_f[1] & input_e[0];
  assign cgp_core_035 = input_a[0] ^ input_e[2];
  assign cgp_core_036 = ~input_e[2];
  assign cgp_core_039 = ~input_f[2];
  assign cgp_core_040 = input_e[2] | input_d[1];
  assign cgp_core_041 = input_e[0] ^ input_d[1];
  assign cgp_core_043 = input_c[2] | cgp_core_039;
  assign cgp_core_044 = input_a[2] | cgp_core_043;
  assign cgp_core_045 = input_a[2] & cgp_core_043;
  assign cgp_core_046 = ~(input_c[0] ^ input_f[1]);
  assign cgp_core_047 = ~(input_f[1] & input_f[2]);
  assign cgp_core_048_not = ~input_e[2];
  assign cgp_core_051 = ~(input_d[2] ^ input_d[2]);
  assign cgp_core_052 = ~(input_b[2] ^ input_a[2]);
  assign cgp_core_053_not = ~input_c[0];
  assign cgp_core_055 = input_d[0] & input_e[2];
  assign cgp_core_056 = ~(input_f[1] ^ input_c[0]);
  assign cgp_core_057 = ~(input_d[0] | input_c[1]);
  assign cgp_core_058 = input_c[0] ^ input_d[2];
  assign cgp_core_060 = ~(input_c[0] & input_e[2]);
  assign cgp_core_063 = input_c[2] ^ input_e[0];
  assign cgp_core_064 = input_d[1] | input_a[2];
  assign cgp_core_065 = ~input_c[0];
  assign cgp_core_067 = input_e[0] ^ input_a[0];
  assign cgp_core_068 = ~input_a[1];
  assign cgp_core_069 = ~(input_d[2] ^ input_b[2]);
  assign cgp_core_070 = ~(input_b[0] ^ input_c[2]);
  assign cgp_core_071 = input_d[2] & input_b[2];
  assign cgp_core_072 = ~cgp_core_071;
  assign cgp_core_073 = cgp_core_045 & cgp_core_072;
  assign cgp_core_074 = ~(cgp_core_045 ^ cgp_core_071);
  assign cgp_core_075 = ~(input_e[0] ^ input_b[0]);
  assign cgp_core_076 = cgp_core_044 & input_e[2];
  assign cgp_core_077 = cgp_core_076 & cgp_core_074;
  assign cgp_core_078 = ~input_e[0];
  assign cgp_core_079 = ~(input_c[1] | input_a[2]);
  assign cgp_core_080 = ~input_f[0];
  assign cgp_core_082 = ~(input_e[1] & input_b[2]);
  assign cgp_core_084 = ~(input_b[1] ^ input_d[1]);
  assign cgp_core_085 = ~input_d[1];
  assign cgp_core_087 = input_e[0] | input_f[2];
  assign cgp_core_088 = ~input_a[1];
  assign cgp_core_089 = ~input_e[0];
  assign cgp_core_090 = input_e[2] ^ input_e[2];
  assign cgp_core_091 = input_b[1] | input_a[0];
  assign cgp_core_092 = input_b[2] | input_e[1];
  assign cgp_core_094 = ~(input_a[2] & input_b[0]);
  assign cgp_core_095 = input_c[0] | input_f[0];
  assign cgp_core_098 = cgp_core_077 | cgp_core_073;
  assign cgp_core_099 = input_d[0] | input_d[2];

  assign cgp_out[0] = cgp_core_098;
endmodule