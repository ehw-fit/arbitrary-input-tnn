module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_069_not;
  wire cgp_core_071;
  wire cgp_core_076;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_088;
  wire cgp_core_095;

  assign cgp_core_019 = ~(input_d[0] | input_h[0]);
  assign cgp_core_020 = input_d[1] ^ input_f[0];
  assign cgp_core_021 = input_f[0] & input_d[1];
  assign cgp_core_022 = ~(input_g[0] & cgp_core_019);
  assign cgp_core_023 = ~(cgp_core_020 & cgp_core_019);
  assign cgp_core_024 = cgp_core_021 | input_g[1];
  assign cgp_core_025 = ~(input_a[0] & input_a[0]);
  assign cgp_core_026 = ~(input_a[0] & input_d[0]);
  assign cgp_core_028 = input_a[1] & cgp_core_022;
  assign cgp_core_031 = input_f[1] | input_d[1];
  assign cgp_core_032 = cgp_core_024 ^ cgp_core_031;
  assign cgp_core_033 = input_g[0] & cgp_core_031;
  assign cgp_core_035 = input_g[0] & input_c[0];
  assign cgp_core_036 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_038 = cgp_core_036 ^ cgp_core_035;
  assign cgp_core_039 = input_h[0] & input_a[1];
  assign cgp_core_041 = input_e[0] ^ input_f[0];
  assign cgp_core_043 = input_f[1] & input_g[1];
  assign cgp_core_044 = input_f[1] & input_g[1];
  assign cgp_core_045 = cgp_core_043 ^ input_f[0];
  assign cgp_core_046 = input_h[1] & input_e[1];
  assign cgp_core_047 = ~(cgp_core_044 | cgp_core_046);
  assign cgp_core_048_not = ~input_e[0];
  assign cgp_core_049 = input_e[0] & cgp_core_041;
  assign cgp_core_050 = input_e[1] ^ cgp_core_045;
  assign cgp_core_051 = input_h[0] & input_g[1];
  assign cgp_core_052 = input_b[0] ^ cgp_core_049;
  assign cgp_core_056 = input_a[0] & input_e[1];
  assign cgp_core_057 = ~(input_h[1] ^ cgp_core_048_not);
  assign cgp_core_059 = cgp_core_038 ^ cgp_core_052;
  assign cgp_core_060 = cgp_core_038 & cgp_core_052;
  assign cgp_core_069_not = ~cgp_core_056;
  assign cgp_core_071 = ~input_c[1];
  assign cgp_core_076 = ~(input_e[0] & cgp_core_069_not);
  assign cgp_core_083 = ~input_d[1];
  assign cgp_core_084 = ~(input_b[0] ^ cgp_core_083);
  assign cgp_core_088 = ~input_h[1];
  assign cgp_core_095 = input_a[0] | input_g[1];

  assign cgp_out[0] = 1'b0;
endmodule