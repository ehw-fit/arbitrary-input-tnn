module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044_not;
  wire cgp_core_045_not;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063_not;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_019 = ~(input_c[1] ^ input_c[1]);
  assign cgp_core_020 = ~(input_d[1] & input_c[1]);
  assign cgp_core_021 = ~(input_g[0] | input_b[1]);
  assign cgp_core_022 = input_e[0] ^ cgp_core_021;
  assign cgp_core_026 = ~(input_a[1] ^ input_d[0]);
  assign cgp_core_027 = input_c[1] ^ input_c[1];
  assign cgp_core_029 = ~(input_a[1] | input_a[0]);
  assign cgp_core_033 = ~(input_g[1] & cgp_core_027);
  assign cgp_core_034 = input_a[0] ^ input_d[1];
  assign cgp_core_035 = ~(input_b[1] | input_c[1]);
  assign cgp_core_037 = ~(input_e[0] | input_e[0]);
  assign cgp_core_038 = cgp_core_022 & input_c[0];
  assign cgp_core_039 = ~input_d[0];
  assign cgp_core_041 = ~(input_a[0] | input_d[1]);
  assign cgp_core_043 = ~(input_f[1] | input_c[1]);
  assign cgp_core_044_not = ~input_c[0];
  assign cgp_core_045_not = ~input_g[0];
  assign cgp_core_046 = ~(input_f[1] | input_b[0]);
  assign cgp_core_047 = input_d[1] ^ input_b[1];
  assign cgp_core_049 = ~(input_f[1] | input_a[0]);
  assign cgp_core_052 = input_e[1] & input_e[0];
  assign cgp_core_057 = input_c[1] | input_g[1];
  assign cgp_core_058 = ~input_d[1];
  assign cgp_core_059 = ~input_d[1];
  assign cgp_core_060 = ~(input_f[1] ^ input_c[1]);
  assign cgp_core_062 = input_f[1] & input_e[1];
  assign cgp_core_063_not = ~cgp_core_062;
  assign cgp_core_064 = cgp_core_039 & input_b[1];
  assign cgp_core_067 = input_d[1] & input_f[1];
  assign cgp_core_068 = ~(cgp_core_067 ^ input_a[0]);
  assign cgp_core_069 = ~input_f[1];
  assign cgp_core_071 = input_b[1] & input_b[0];
  assign cgp_core_075 = ~input_f[0];
  assign cgp_core_076 = input_c[1] | input_a[1];
  assign cgp_core_077 = ~(input_b[0] & input_f[1]);
  assign cgp_core_079 = ~(input_g[0] & input_g[0]);

  assign cgp_out[0] = 1'b1;
endmodule