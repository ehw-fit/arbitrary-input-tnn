module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_038_not;
  wire cgp_core_042;

  assign cgp_core_014 = input_a[0] & input_b[0];
  assign cgp_core_015 = ~(input_a[1] | input_b[1]);
  assign cgp_core_016 = input_c[1] & input_b[0];
  assign cgp_core_017 = cgp_core_014 | cgp_core_016;
  assign cgp_core_018 = input_a[2] | input_c[2];
  assign cgp_core_019 = input_a[2] & input_c[2];
  assign cgp_core_020 = cgp_core_018 | cgp_core_017;
  assign cgp_core_021 = cgp_core_018 & cgp_core_017;
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_023 = ~(input_a[2] & input_c[0]);
  assign cgp_core_024 = ~cgp_core_022;
  assign cgp_core_025 = ~cgp_core_020;
  assign cgp_core_026 = input_b[2] & cgp_core_025;
  assign cgp_core_028 = ~(input_b[2] ^ cgp_core_020);
  assign cgp_core_029 = cgp_core_028 & cgp_core_024;
  assign cgp_core_031 = input_b[0] ^ input_a[0];
  assign cgp_core_032 = input_b[0] & cgp_core_029;
  assign cgp_core_033 = input_c[1] & input_c[2];
  assign cgp_core_034 = input_b[0] | input_a[2];
  assign cgp_core_038_not = ~input_c[2];
  assign cgp_core_042 = cgp_core_032 | cgp_core_026;

  assign cgp_out[0] = cgp_core_042;
endmodule