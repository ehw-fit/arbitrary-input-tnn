module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021_not;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_060_not;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067_not;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_076;
  wire cgp_core_079;
  wire cgp_core_083;

  assign cgp_core_016 = ~input_f[0];
  assign cgp_core_017 = ~(input_f[0] ^ input_g[0]);
  assign cgp_core_019 = ~(input_e[1] & input_f[0]);
  assign cgp_core_020 = ~input_f[0];
  assign cgp_core_021_not = ~input_a[1];
  assign cgp_core_022 = input_b[1] | input_b[1];
  assign cgp_core_023 = ~(input_e[1] & input_b[0]);
  assign cgp_core_025 = ~input_c[1];
  assign cgp_core_027 = ~(input_b[1] ^ input_f[1]);
  assign cgp_core_028 = input_e[0] ^ input_b[0];
  assign cgp_core_029 = input_e[1] | input_c[0];
  assign cgp_core_030 = input_a[1] & input_a[0];
  assign cgp_core_031 = ~input_e[1];
  assign cgp_core_032 = ~(input_b[1] & input_e[0]);
  assign cgp_core_034 = input_e[1] & input_g[0];
  assign cgp_core_035 = input_c[0] & input_e[0];
  assign cgp_core_036 = input_g[1] | input_c[1];
  assign cgp_core_037 = input_c[0] | cgp_core_036;
  assign cgp_core_038 = cgp_core_029 & cgp_core_036;
  assign cgp_core_039 = ~(input_d[0] & input_e[0]);
  assign cgp_core_040 = ~(input_f[1] | input_c[0]);
  assign cgp_core_041 = input_c[1] ^ input_e[1];
  assign cgp_core_042 = ~input_f[1];
  assign cgp_core_043_not = ~input_e[1];
  assign cgp_core_044 = ~(input_g[0] & input_e[1]);
  assign cgp_core_045 = input_a[1] | input_d[1];
  assign cgp_core_046 = input_e[1] | cgp_core_037;
  assign cgp_core_048 = cgp_core_046 | cgp_core_045;
  assign cgp_core_049 = cgp_core_046 & cgp_core_045;
  assign cgp_core_051 = cgp_core_038 | cgp_core_049;
  assign cgp_core_052 = input_b[1] & input_g[1];
  assign cgp_core_053 = ~(input_f[1] ^ input_f[1]);
  assign cgp_core_054 = input_f[0] ^ input_d[1];
  assign cgp_core_056 = input_b[1] & input_f[1];
  assign cgp_core_060_not = ~input_g[1];
  assign cgp_core_062 = ~(input_e[1] & input_b[0]);
  assign cgp_core_063 = input_d[0] & input_a[1];
  assign cgp_core_064 = ~cgp_core_056;
  assign cgp_core_065 = cgp_core_048 & cgp_core_064;
  assign cgp_core_067_not = ~input_g[1];
  assign cgp_core_068 = ~input_f[0];
  assign cgp_core_069 = ~(input_d[0] & input_f[0]);
  assign cgp_core_070 = input_g[0] & input_a[0];
  assign cgp_core_071 = cgp_core_070 & input_d[0];
  assign cgp_core_073 = ~(input_e[0] & input_d[0]);
  assign cgp_core_074_not = ~input_c[0];
  assign cgp_core_076 = ~(input_g[0] ^ input_f[1]);
  assign cgp_core_079 = cgp_core_071 | cgp_core_065;
  assign cgp_core_083 = cgp_core_079 | cgp_core_051;

  assign cgp_out[0] = cgp_core_083;
endmodule