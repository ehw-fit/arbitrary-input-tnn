module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;

  assign cgp_core_016 = input_a[1] | input_a[2];
  assign cgp_core_017 = input_a[1] & input_a[2];
  assign cgp_core_018 = input_a[9] & input_a[3];
  assign cgp_core_019 = input_a[0] & cgp_core_016;
  assign cgp_core_020 = cgp_core_017 | cgp_core_019;
  assign cgp_core_023 = input_a[9] & input_a[4];
  assign cgp_core_024 = input_a[5] ^ input_a[6];
  assign cgp_core_025 = input_a[5] & input_a[6];
  assign cgp_core_028 = cgp_core_023 ^ cgp_core_025;
  assign cgp_core_029 = cgp_core_023 & cgp_core_025;
  assign cgp_core_031 = input_a[10] & input_a[7];
  assign cgp_core_034 = input_a[11] & cgp_core_024;
  assign cgp_core_035 = cgp_core_020 ^ cgp_core_028;
  assign cgp_core_036 = cgp_core_020 & cgp_core_028;
  assign cgp_core_037 = cgp_core_035 ^ cgp_core_034;
  assign cgp_core_038 = cgp_core_035 & cgp_core_034;
  assign cgp_core_039 = cgp_core_036 | cgp_core_038;
  assign cgp_core_042 = cgp_core_029 | cgp_core_039;
  assign cgp_core_044 = input_a[6] | input_a[2];
  assign cgp_core_046 = input_a[1] | input_a[7];
  assign cgp_core_047 = ~input_a[2];
  assign cgp_core_048 = input_a[12] | input_a[11];
  assign cgp_core_051 = input_a[2] & input_a[8];
  assign cgp_core_052 = input_a[10] & input_a[7];
  assign cgp_core_053 = input_a[12] & input_a[9];
  assign cgp_core_054 = ~input_a[9];
  assign cgp_core_055 = ~input_a[13];
  assign cgp_core_057 = cgp_core_052 ^ input_a[12];
  assign cgp_core_062 = ~(input_a[5] ^ input_a[9]);
  assign cgp_core_063 = ~(input_a[12] | cgp_core_055);
  assign cgp_core_064_not = ~cgp_core_057;
  assign cgp_core_066 = cgp_core_064_not ^ cgp_core_063;
  assign cgp_core_067 = ~(input_a[10] | input_a[3]);
  assign cgp_core_069 = input_a[13] | cgp_core_052;
  assign cgp_core_070 = ~(input_a[10] | input_a[2]);
  assign cgp_core_071 = cgp_core_069 | input_a[12];
  assign cgp_core_073 = ~(input_a[6] | input_a[1]);
  assign cgp_core_075 = input_a[3] & input_a[8];
  assign cgp_core_076 = cgp_core_037 ^ cgp_core_066;
  assign cgp_core_077 = cgp_core_037 & cgp_core_066;
  assign cgp_core_078 = cgp_core_076 ^ cgp_core_075;
  assign cgp_core_079 = cgp_core_076 & cgp_core_075;
  assign cgp_core_080 = cgp_core_077 | cgp_core_079;
  assign cgp_core_081 = cgp_core_042 ^ cgp_core_071;
  assign cgp_core_082 = cgp_core_042 & cgp_core_071;
  assign cgp_core_083 = cgp_core_081 ^ cgp_core_080;
  assign cgp_core_084 = cgp_core_081 & cgp_core_080;
  assign cgp_core_085 = cgp_core_082 | cgp_core_084;
  assign cgp_core_086 = ~input_a[12];

  assign cgp_out[0] = 1'b0;
  assign cgp_out[1] = cgp_core_078;
  assign cgp_out[2] = cgp_core_083;
  assign cgp_out[3] = cgp_core_085;
endmodule