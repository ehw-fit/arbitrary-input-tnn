module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_030;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_016 = input_d[0] ^ input_g[1];
  assign cgp_core_018 = input_c[1] ^ input_e[1];
  assign cgp_core_019 = input_c[1] & input_e[1];
  assign cgp_core_025 = input_a[1] ^ cgp_core_018;
  assign cgp_core_026 = input_a[1] & cgp_core_018;
  assign cgp_core_030 = cgp_core_019 | cgp_core_026;
  assign cgp_core_032_not = ~input_b[1];
  assign cgp_core_033 = ~(input_a[0] | input_g[0]);
  assign cgp_core_034 = input_g[1] | input_e[0];
  assign cgp_core_035 = input_b[1] & input_g[0];
  assign cgp_core_037 = ~input_a[0];
  assign cgp_core_040 = ~(input_g[0] & input_f[1]);
  assign cgp_core_041 = input_f[1] | input_g[1];
  assign cgp_core_042 = input_f[1] & input_g[1];
  assign cgp_core_043 = input_d[1] ^ input_e[0];
  assign cgp_core_044 = cgp_core_041 & input_d[1];
  assign cgp_core_045 = cgp_core_042 | cgp_core_044;
  assign cgp_core_046 = ~(input_e[0] & input_e[0]);
  assign cgp_core_047 = input_b[0] | input_e[0];
  assign cgp_core_048 = input_g[1] | input_c[1];
  assign cgp_core_050 = ~(input_g[0] ^ input_e[0]);
  assign cgp_core_051 = ~(input_f[0] ^ input_d[0]);
  assign cgp_core_053 = cgp_core_035 | cgp_core_045;
  assign cgp_core_057 = ~input_e[1];
  assign cgp_core_058 = ~(input_a[1] | input_a[0]);
  assign cgp_core_059 = input_f[0] ^ input_c[1];
  assign cgp_core_061 = ~cgp_core_053;
  assign cgp_core_062 = cgp_core_030 & cgp_core_061;
  assign cgp_core_068 = cgp_core_025 & cgp_core_030;
  assign cgp_core_070 = input_b[0] | input_a[0];
  assign cgp_core_071 = ~(input_f[1] ^ input_a[0]);
  assign cgp_core_073 = ~(input_a[1] | input_g[0]);
  assign cgp_core_077 = ~(input_c[1] ^ input_b[1]);
  assign cgp_core_079 = cgp_core_068 | cgp_core_062;

  assign cgp_out[0] = cgp_core_079;
endmodule