module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017_not = ~input_b[0];
  assign cgp_core_018 = input_a[0] & input_c[2];
  assign cgp_core_019 = input_e[2] ^ input_b[1];
  assign cgp_core_020 = ~(input_a[1] & input_b[1]);
  assign cgp_core_022 = input_b[0] & cgp_core_018;
  assign cgp_core_023 = ~(input_d[0] & input_d[0]);
  assign cgp_core_024 = input_b[1] ^ input_c[2];
  assign cgp_core_027 = input_e[2] & cgp_core_023;
  assign cgp_core_029 = ~(input_d[0] ^ input_e[0]);
  assign cgp_core_030 = input_d[0] & input_c[1];
  assign cgp_core_031 = input_b[2] ^ input_e[1];
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_034 = ~input_b[1];
  assign cgp_core_036 = ~(input_a[0] & input_a[2]);
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038_not = ~cgp_core_036;
  assign cgp_core_040 = input_a[2] | input_d[2];
  assign cgp_core_041 = input_c[0] ^ input_e[1];
  assign cgp_core_042 = input_c[0] & cgp_core_029;
  assign cgp_core_043_not = ~input_e[1];
  assign cgp_core_045 = ~(input_b[2] | input_e[1]);
  assign cgp_core_046 = input_c[2] & input_a[2];
  assign cgp_core_047 = input_d[2] | input_b[2];
  assign cgp_core_048 = input_b[2] ^ input_b[0];
  assign cgp_core_049 = input_c[2] | cgp_core_038_not;
  assign cgp_core_051 = ~cgp_core_048;
  assign cgp_core_053 = input_c[2] ^ input_c[1];
  assign cgp_core_054 = input_b[1] & input_c[1];
  assign cgp_core_055 = ~input_c[0];
  assign cgp_core_056 = ~(input_c[0] & cgp_core_054);
  assign cgp_core_057 = cgp_core_053 ^ input_a[1];
  assign cgp_core_059 = cgp_core_057 & input_e[2];
  assign cgp_core_060 = ~(input_e[0] ^ input_d[2]);
  assign cgp_core_061 = cgp_core_060 & cgp_core_056;
  assign cgp_core_064 = input_c[1] & input_e[0];
  assign cgp_core_065 = ~(input_e[2] ^ input_a[2]);
  assign cgp_core_067 = ~cgp_core_045;
  assign cgp_core_072 = ~(cgp_core_041 | cgp_core_041);
  assign cgp_core_073 = ~(cgp_core_017_not | input_c[2]);
  assign cgp_core_075 = ~(input_c[1] ^ input_e[0]);
  assign cgp_core_079 = input_d[0] | input_c[1];
  assign cgp_core_080 = input_e[1] | input_c[0];

  assign cgp_out[0] = 1'b0;
endmodule