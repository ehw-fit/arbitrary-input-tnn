module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_048_not;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = ~input_g[1];
  assign cgp_core_017 = ~(input_g[0] | input_g[0]);
  assign cgp_core_018 = ~(input_f[0] & input_c[0]);
  assign cgp_core_020 = ~input_b[1];
  assign cgp_core_021 = input_g[0] | input_d[0];
  assign cgp_core_022 = ~(input_e[0] | input_c[0]);
  assign cgp_core_024 = input_a[0] & input_g[1];
  assign cgp_core_028 = input_f[0] ^ input_b[1];
  assign cgp_core_030 = input_c[1] & input_b[1];
  assign cgp_core_031 = ~input_f[0];
  assign cgp_core_032 = input_g[0] | input_e[0];
  assign cgp_core_034 = ~(input_d[1] ^ input_a[1]);
  assign cgp_core_036 = ~(input_d[0] ^ input_d[1]);
  assign cgp_core_037 = ~(input_e[1] & input_a[1]);
  assign cgp_core_038 = ~(input_g[0] & input_e[1]);
  assign cgp_core_039 = ~(input_c[1] | input_e[1]);
  assign cgp_core_041 = ~input_a[0];
  assign cgp_core_043 = ~(input_a[0] ^ input_e[0]);
  assign cgp_core_046 = input_g[0] | input_d[0];
  assign cgp_core_048_not = ~input_f[1];
  assign cgp_core_054_not = ~input_d[1];
  assign cgp_core_055 = ~input_c[0];
  assign cgp_core_056 = ~(input_d[0] ^ input_d[1]);
  assign cgp_core_057 = ~input_b[0];
  assign cgp_core_058 = ~input_a[0];
  assign cgp_core_059 = input_e[1] & input_f[0];
  assign cgp_core_060 = input_b[1] ^ input_c[0];
  assign cgp_core_061 = ~(input_e[1] ^ input_a[0]);
  assign cgp_core_063 = input_b[0] | input_d[0];
  assign cgp_core_064 = input_d[0] & input_f[0];
  assign cgp_core_065 = input_c[0] & input_b[1];
  assign cgp_core_067 = input_e[1] | input_b[1];
  assign cgp_core_068 = input_f[0] | input_a[1];
  assign cgp_core_069 = input_f[1] | input_d[0];
  assign cgp_core_070 = ~input_f[0];
  assign cgp_core_073 = input_d[0] ^ input_a[1];
  assign cgp_core_074_not = ~input_b[0];
  assign cgp_core_076 = ~(input_c[1] | input_a[1]);
  assign cgp_core_077 = ~input_c[0];
  assign cgp_core_078 = input_c[1] | input_g[1];
  assign cgp_core_079 = input_e[1] | cgp_core_078;

  assign cgp_out[0] = cgp_core_079;
endmodule