parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 12,
parameter FEAT_BITS = 3,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1470
