module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_055_not;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_087;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_095;
  wire cgp_core_096;

  assign cgp_core_018 = input_d[1] & input_f[0];
  assign cgp_core_019 = ~input_b[1];
  assign cgp_core_020 = ~input_c[0];
  assign cgp_core_021 = input_h[0] ^ input_f[1];
  assign cgp_core_022 = ~(input_d[1] & input_h[1]);
  assign cgp_core_024 = input_e[0] | input_e[1];
  assign cgp_core_025 = input_e[1] | input_g[1];
  assign cgp_core_026 = ~(input_c[1] ^ input_f[0]);
  assign cgp_core_027 = input_d[0] | input_d[1];
  assign cgp_core_028 = input_b[1] & input_a[0];
  assign cgp_core_029 = input_e[0] & input_d[0];
  assign cgp_core_030 = input_h[1] & input_g[0];
  assign cgp_core_031 = ~(input_d[1] | input_c[1]);
  assign cgp_core_032 = input_a[0] & input_g[0];
  assign cgp_core_034 = input_a[0] & input_d[0];
  assign cgp_core_039 = input_g[0] ^ input_e[1];
  assign cgp_core_040 = ~(input_h[0] | input_b[0]);
  assign cgp_core_042 = input_h[0] | input_b[1];
  assign cgp_core_043 = input_f[1] | input_g[1];
  assign cgp_core_044 = input_f[1] & input_g[1];
  assign cgp_core_045 = ~(input_a[1] & input_d[1]);
  assign cgp_core_046 = cgp_core_043 & input_c[1];
  assign cgp_core_047 = cgp_core_044 | cgp_core_046;
  assign cgp_core_049 = ~input_c[1];
  assign cgp_core_050_not = ~input_b[1];
  assign cgp_core_051 = ~(input_b[0] & input_h[1]);
  assign cgp_core_053 = ~(input_e[0] & input_b[1]);
  assign cgp_core_055_not = ~input_e[0];
  assign cgp_core_057 = ~(input_a[1] ^ input_f[0]);
  assign cgp_core_058 = ~input_d[0];
  assign cgp_core_060 = input_b[0] | input_c[0];
  assign cgp_core_061 = input_e[0] ^ input_d[1];
  assign cgp_core_062 = ~(input_d[1] | input_e[1]);
  assign cgp_core_067 = input_b[1] & input_e[1];
  assign cgp_core_069 = cgp_core_047 | cgp_core_067;
  assign cgp_core_070 = ~(input_e[1] & input_d[0]);
  assign cgp_core_073 = ~cgp_core_069;
  assign cgp_core_074 = input_h[1] & cgp_core_073;
  assign cgp_core_075 = cgp_core_074 & input_d[1];
  assign cgp_core_076 = input_d[0] | input_a[0];
  assign cgp_core_077 = ~(input_e[0] | input_c[0]);
  assign cgp_core_078 = input_b[0] ^ input_e[1];
  assign cgp_core_081 = input_d[1] & input_f[1];
  assign cgp_core_082 = input_a[1] & input_f[0];
  assign cgp_core_084 = input_b[1] | input_b[0];
  assign cgp_core_087 = input_f[1] & input_c[1];
  assign cgp_core_092 = input_g[0] & input_c[0];
  assign cgp_core_093 = input_b[0] & input_b[0];
  assign cgp_core_095 = ~input_e[1];
  assign cgp_core_096 = ~(input_f[1] | input_d[0]);

  assign cgp_out[0] = cgp_core_075;
endmodule