module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_014 = ~(input_a[0] ^ input_b[1]);
  assign cgp_core_015 = ~(input_a[0] | input_a[0]);
  assign cgp_core_016 = ~(input_b[1] & input_b[1]);
  assign cgp_core_018 = ~(input_d[2] & input_b[1]);
  assign cgp_core_020 = ~(input_c[2] & input_a[2]);
  assign cgp_core_021 = ~input_c[1];
  assign cgp_core_022 = ~(input_d[1] ^ input_d[0]);
  assign cgp_core_023 = ~(input_d[2] | input_a[2]);
  assign cgp_core_024 = input_a[2] & input_b[1];
  assign cgp_core_025 = input_b[2] | cgp_core_024;
  assign cgp_core_026 = input_c[2] ^ input_a[1];
  assign cgp_core_028 = ~(input_d[1] & input_c[0]);
  assign cgp_core_029 = input_d[2] | input_a[0];
  assign cgp_core_030 = input_c[0] ^ input_b[2];
  assign cgp_core_031 = ~(input_c[0] ^ input_b[2]);
  assign cgp_core_033 = ~(input_a[0] & input_d[2]);
  assign cgp_core_034 = ~(input_a[0] ^ input_b[0]);
  assign cgp_core_036 = ~(input_a[0] ^ input_b[0]);
  assign cgp_core_038 = ~input_c[2];
  assign cgp_core_039 = cgp_core_025 & cgp_core_038;
  assign cgp_core_040 = ~(cgp_core_025 ^ input_c[2]);
  assign cgp_core_041 = ~input_d[2];
  assign cgp_core_043 = cgp_core_041 & cgp_core_040;
  assign cgp_core_045 = input_a[2] | input_d[2];
  assign cgp_core_046 = input_a[1] & input_b[1];
  assign cgp_core_047 = ~(input_b[1] & input_d[0]);
  assign cgp_core_050_not = ~input_d[2];
  assign cgp_core_051 = ~(input_b[1] & input_c[1]);
  assign cgp_core_058 = cgp_core_043 | cgp_core_039;
  assign cgp_core_059 = ~(input_c[2] | input_c[1]);

  assign cgp_out[0] = cgp_core_058;
endmodule