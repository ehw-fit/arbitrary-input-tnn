module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_012;
  wire cgp_core_014;
  wire cgp_core_018;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_054_not;

  assign cgp_core_012 = ~input_b[0];
  assign cgp_core_014 = input_c[0] & input_a[0];
  assign cgp_core_018 = input_c[0] | input_a[0];
  assign cgp_core_023_not = ~input_d[0];
  assign cgp_core_024 = ~(input_c[1] | input_c[0]);
  assign cgp_core_026 = ~(input_d[1] | input_e[1]);
  assign cgp_core_027 = ~(input_b[0] ^ input_a[0]);
  assign cgp_core_030 = ~(input_d[1] & input_e[1]);
  assign cgp_core_031 = input_e[1] ^ input_a[0];
  assign cgp_core_032 = ~(input_e[0] | input_c[0]);
  assign cgp_core_034 = input_c[0] & input_b[0];
  assign cgp_core_037 = ~input_c[1];
  assign cgp_core_038 = input_c[0] & input_b[1];
  assign cgp_core_039 = input_c[1] ^ input_a[0];
  assign cgp_core_040 = ~(input_d[1] & input_c[1]);
  assign cgp_core_042 = ~input_c[1];
  assign cgp_core_043 = input_e[0] & input_b[0];
  assign cgp_core_045 = ~(input_b[0] & input_d[1]);
  assign cgp_core_046 = ~input_d[0];
  assign cgp_core_048 = input_d[1] ^ input_e[0];
  assign cgp_core_049 = input_d[0] & input_c[1];
  assign cgp_core_050 = ~(cgp_core_012 & input_b[0]);
  assign cgp_core_054_not = ~input_d[1];

  assign cgp_out[0] = 1'b0;
endmodule