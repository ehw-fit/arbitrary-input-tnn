module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_018_not;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_029;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045_not;
  wire cgp_core_047;
  wire cgp_core_048_not;
  wire cgp_core_049;
  wire cgp_core_051_not;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_059;

  assign cgp_core_014 = ~input_b[1];
  assign cgp_core_016_not = ~input_a[1];
  assign cgp_core_017 = input_b[0] ^ input_a[1];
  assign cgp_core_018_not = ~input_c[0];
  assign cgp_core_019 = input_c[1] | input_c[2];
  assign cgp_core_020 = input_c[2] & input_d[2];
  assign cgp_core_021 = ~(input_b[0] & input_c[1]);
  assign cgp_core_023 = input_a[2] | input_b[1];
  assign cgp_core_024 = ~(input_b[0] ^ input_a[2]);
  assign cgp_core_026 = ~(input_d[2] & input_b[2]);
  assign cgp_core_027_not = ~input_d[0];
  assign cgp_core_029 = input_b[1] & input_d[0];
  assign cgp_core_033 = input_a[1] & input_a[2];
  assign cgp_core_034 = ~(input_b[2] ^ input_c[0]);
  assign cgp_core_035 = ~(input_d[1] & input_b[1]);
  assign cgp_core_036 = input_b[0] ^ input_a[0];
  assign cgp_core_037 = ~input_b[0];
  assign cgp_core_040 = input_c[0] & input_b[1];
  assign cgp_core_042 = ~input_c[2];
  assign cgp_core_043 = ~(input_c[2] | input_d[2]);
  assign cgp_core_045_not = ~input_c[0];
  assign cgp_core_047 = ~(input_d[2] ^ input_a[0]);
  assign cgp_core_048_not = ~input_d[0];
  assign cgp_core_049 = input_b[1] & input_a[1];
  assign cgp_core_051_not = ~input_a[2];
  assign cgp_core_052 = ~(input_d[1] ^ input_a[0]);
  assign cgp_core_053 = ~(input_c[0] | input_a[0]);
  assign cgp_core_054 = ~input_a[1];
  assign cgp_core_057 = ~(input_b[0] | input_b[0]);
  assign cgp_core_059 = input_b[2] | cgp_core_043;

  assign cgp_out[0] = cgp_core_059;
endmodule