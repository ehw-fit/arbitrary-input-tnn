module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_020_not;
  wire cgp_core_022_not;
  wire cgp_core_024_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_015 = ~input_a[0];
  assign cgp_core_016 = input_a[1] & input_a[9];
  assign cgp_core_018 = input_a[5] & input_a[3];
  assign cgp_core_020_not = ~input_a[10];
  assign cgp_core_022_not = ~input_a[4];
  assign cgp_core_024_not = ~input_a[1];
  assign cgp_core_028 = ~(input_a[6] | input_a[1]);
  assign cgp_core_029 = input_a[6] | input_a[0];
  assign cgp_core_032 = ~input_a[4];
  assign cgp_core_033 = input_a[1] & input_a[3];
  assign cgp_core_034 = input_a[1] & input_a[2];
  assign cgp_core_035 = input_a[6] ^ input_a[5];
  assign cgp_core_037 = ~input_a[5];
  assign cgp_core_039 = input_a[11] & input_a[0];
  assign cgp_core_040 = input_a[0] | input_a[11];
  assign cgp_core_041 = ~(input_a[5] | input_a[11]);
  assign cgp_core_042_not = ~input_a[7];
  assign cgp_core_044 = input_a[8] ^ input_a[2];
  assign cgp_core_045 = input_a[0] ^ input_a[0];
  assign cgp_core_046 = ~(input_a[2] ^ input_a[6]);
  assign cgp_core_047 = ~(input_a[9] ^ input_a[5]);
  assign cgp_core_048 = input_a[2] & input_a[4];
  assign cgp_core_049 = input_a[6] & input_a[8];
  assign cgp_core_050 = ~(input_a[2] | input_a[10]);
  assign cgp_core_052 = ~input_a[2];
  assign cgp_core_055 = input_a[1] ^ input_a[6];
  assign cgp_core_056 = input_a[0] | input_a[3];
  assign cgp_core_058 = input_a[6] | input_a[11];
  assign cgp_core_061 = input_a[4] & input_a[0];
  assign cgp_core_063 = ~(input_a[3] & input_a[1]);
  assign cgp_core_067 = ~(input_a[10] & input_a[3]);
  assign cgp_core_070 = ~(input_a[1] ^ input_a[0]);
  assign cgp_core_071 = input_a[9] ^ input_a[1];
  assign cgp_core_074 = input_a[2] ^ input_a[5];
  assign cgp_core_075 = input_a[6] & input_a[10];
  assign cgp_core_076 = ~(input_a[7] ^ input_a[1]);
  assign cgp_core_077 = ~input_a[5];
  assign cgp_core_078 = input_a[3] & input_a[11];

  assign cgp_out[0] = 1'b0;
  assign cgp_out[1] = input_a[10];
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = 1'b0;
endmodule