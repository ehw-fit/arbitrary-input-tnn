module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_058_not;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_081;
  wire cgp_core_082_not;
  wire cgp_core_083;
  wire cgp_core_084_not;
  wire cgp_core_085_not;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_095;

  assign cgp_core_020 = ~(input_a[0] | input_b[0]);
  assign cgp_core_022 = ~(input_b[0] | input_b[0]);
  assign cgp_core_023 = ~input_a[2];
  assign cgp_core_025 = ~input_a[2];
  assign cgp_core_027 = input_d[0] ^ input_c[0];
  assign cgp_core_029 = input_a[0] & input_a[0];
  assign cgp_core_030 = input_d[1] | input_a[1];
  assign cgp_core_031 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_033 = input_e[2] & input_d[0];
  assign cgp_core_034 = ~(input_c[1] & input_a[0]);
  assign cgp_core_035 = input_d[2] & input_e[2];
  assign cgp_core_037 = ~(cgp_core_034 ^ cgp_core_033);
  assign cgp_core_039 = input_c[2] & input_f[2];
  assign cgp_core_041 = input_d[2] | input_b[2];
  assign cgp_core_042 = input_a[0] & input_b[0];
  assign cgp_core_045 = ~input_a[0];
  assign cgp_core_049 = ~(input_f[1] ^ input_b[1]);
  assign cgp_core_051 = input_e[0] & input_f[2];
  assign cgp_core_052 = ~(input_e[2] | input_e[0]);
  assign cgp_core_055 = ~(cgp_core_052 & input_f[0]);
  assign cgp_core_058_not = ~input_d[0];
  assign cgp_core_059 = ~input_f[1];
  assign cgp_core_060 = cgp_core_058_not ^ input_d[2];
  assign cgp_core_061 = ~(cgp_core_058_not | input_c[0]);
  assign cgp_core_062 = input_a[0] ^ input_a[1];
  assign cgp_core_065 = input_d[2] & input_f[1];
  assign cgp_core_066 = input_c[1] & input_b[0];
  assign cgp_core_067 = input_e[0] | input_b[2];
  assign cgp_core_069 = ~(input_c[1] | input_c[0]);
  assign cgp_core_072 = ~(cgp_core_069 ^ input_e[2]);
  assign cgp_core_073 = ~cgp_core_072;
  assign cgp_core_074 = ~input_e[1];
  assign cgp_core_075 = ~input_f[1];
  assign cgp_core_076 = input_e[2] & input_b[1];
  assign cgp_core_081 = cgp_core_029 & input_e[2];
  assign cgp_core_082_not = ~input_a[2];
  assign cgp_core_083 = ~input_a[0];
  assign cgp_core_084_not = ~input_f[2];
  assign cgp_core_085_not = ~input_b[1];
  assign cgp_core_088 = ~(input_e[1] & input_e[1]);
  assign cgp_core_090 = input_e[2] ^ input_c[1];
  assign cgp_core_095 = input_a[1] | cgp_core_082_not;

  assign cgp_out[0] = 1'b0;
endmodule