module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032_not;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067_not;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_078;

  assign cgp_core_017 = ~(input_d[0] | input_e[0]);
  assign cgp_core_019 = input_c[0] & input_b[0];
  assign cgp_core_020 = ~(input_a[0] & input_b[1]);
  assign cgp_core_021 = input_a[0] ^ input_c[1];
  assign cgp_core_023 = ~input_a[0];
  assign cgp_core_024 = input_a[0] & input_d[0];
  assign cgp_core_026 = input_d[0] ^ input_d[0];
  assign cgp_core_028 = input_b[1] & input_g[1];
  assign cgp_core_029 = ~(input_a[0] ^ cgp_core_028);
  assign cgp_core_030 = ~input_f[0];
  assign cgp_core_031 = input_g[1] & cgp_core_029;
  assign cgp_core_032_not = ~input_c[0];
  assign cgp_core_033 = ~input_e[0];
  assign cgp_core_034 = input_f[0] ^ input_d[1];
  assign cgp_core_035 = input_c[0] & input_c[1];
  assign cgp_core_036 = cgp_core_034 & input_c[0];
  assign cgp_core_037 = input_f[0] & input_c[1];
  assign cgp_core_038 = ~(cgp_core_035 | input_b[1]);
  assign cgp_core_039 = ~(input_b[1] | input_e[0]);
  assign cgp_core_040 = input_d[0] & input_g[1];
  assign cgp_core_041 = ~input_f[1];
  assign cgp_core_042 = input_f[1] & input_d[0];
  assign cgp_core_043 = ~(cgp_core_041 & input_g[1]);
  assign cgp_core_044 = input_a[0] & cgp_core_040;
  assign cgp_core_045 = input_e[1] | input_c[0];
  assign cgp_core_049 = ~cgp_core_036;
  assign cgp_core_050 = input_d[0] ^ input_f[0];
  assign cgp_core_052 = input_b[1] & input_a[1];
  assign cgp_core_053 = ~(cgp_core_038 & input_d[1]);
  assign cgp_core_054 = ~(input_a[1] | input_e[1]);
  assign cgp_core_055 = cgp_core_053 ^ cgp_core_052;
  assign cgp_core_056 = ~(input_g[0] | input_g[1]);
  assign cgp_core_057 = cgp_core_054 ^ input_f[1];
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = input_g[1] ^ input_d[0];
  assign cgp_core_060 = input_a[0] & cgp_core_057;
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_063 = ~input_e[1];
  assign cgp_core_064_not = ~cgp_core_055;
  assign cgp_core_065 = input_d[0] & input_c[0];
  assign cgp_core_066 = ~(cgp_core_050 & input_a[1]);
  assign cgp_core_067_not = ~input_a[1];
  assign cgp_core_068 = input_f[0] & cgp_core_065;
  assign cgp_core_069_not = ~cgp_core_050;
  assign cgp_core_070 = input_a[1] & cgp_core_065;
  assign cgp_core_072 = input_d[0] & input_c[0];
  assign cgp_core_073 = input_a[0] ^ cgp_core_070;
  assign cgp_core_078 = ~(cgp_core_063 | input_d[0]);

  assign cgp_out[0] = 1'b0;
endmodule