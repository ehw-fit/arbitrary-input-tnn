module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_080;
  wire cgp_core_083;

  assign cgp_core_018 = ~(input_e[0] ^ input_b[0]);
  assign cgp_core_021 = input_a[1] & input_c[1];
  assign cgp_core_023 = ~(input_e[0] ^ input_e[0]);
  assign cgp_core_024 = input_a[0] & input_g[0];
  assign cgp_core_025 = input_e[1] | input_g[1];
  assign cgp_core_026 = input_e[1] & input_g[1];
  assign cgp_core_027 = cgp_core_025 | cgp_core_024;
  assign cgp_core_028 = cgp_core_025 & input_g[0];
  assign cgp_core_029 = cgp_core_026 | cgp_core_028;
  assign cgp_core_030 = input_c[0] ^ input_c[0];
  assign cgp_core_032 = input_d[1] | cgp_core_027;
  assign cgp_core_033 = input_d[1] & cgp_core_027;
  assign cgp_core_034 = ~input_g[1];
  assign cgp_core_035 = cgp_core_032 & input_e[0];
  assign cgp_core_036 = cgp_core_033 | cgp_core_035;
  assign cgp_core_039 = ~(input_f[0] ^ input_b[1]);
  assign cgp_core_042 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_043 = input_b[1] ^ input_c[0];
  assign cgp_core_045 = ~input_b[0];
  assign cgp_core_046 = cgp_core_021 | cgp_core_036;
  assign cgp_core_047 = input_e[1] ^ input_e[1];
  assign cgp_core_048 = input_c[0] | input_d[0];
  assign cgp_core_051 = cgp_core_029 | cgp_core_046;
  assign cgp_core_052 = ~(input_f[1] | input_b[1]);
  assign cgp_core_054 = input_c[0] ^ input_a[1];
  assign cgp_core_055 = input_b[1] ^ input_f[1];
  assign cgp_core_057 = cgp_core_055 ^ input_c[0];
  assign cgp_core_059 = ~input_e[1];
  assign cgp_core_060 = input_d[1] | input_g[1];
  assign cgp_core_062 = ~input_b[1];
  assign cgp_core_066 = cgp_core_048 & cgp_core_062;
  assign cgp_core_067 = ~(cgp_core_048 ^ input_b[1]);
  assign cgp_core_070 = ~(input_a[1] | input_a[0]);
  assign cgp_core_071 = ~(input_g[0] & input_d[0]);
  assign cgp_core_072 = ~(cgp_core_043 ^ cgp_core_057);
  assign cgp_core_073 = cgp_core_072 & cgp_core_067;
  assign cgp_core_075 = ~(input_f[0] & input_d[0]);
  assign cgp_core_077 = input_b[1] ^ input_g[0];
  assign cgp_core_080 = cgp_core_073 | cgp_core_066;
  assign cgp_core_083 = cgp_core_080 | cgp_core_051;

  assign cgp_out[0] = cgp_core_083;
endmodule