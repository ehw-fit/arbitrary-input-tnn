module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068_not;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_079_not;

  assign cgp_core_017 = input_c[0] & input_d[0];
  assign cgp_core_018 = input_e[0] ^ input_b[1];
  assign cgp_core_022 = input_a[1] | input_e[0];
  assign cgp_core_023 = ~input_b[2];
  assign cgp_core_024_not = ~input_b[2];
  assign cgp_core_025 = input_c[0] | input_b[2];
  assign cgp_core_026 = ~(input_e[0] | input_c[2]);
  assign cgp_core_027 = ~input_c[0];
  assign cgp_core_029 = ~(input_a[1] | input_e[0]);
  assign cgp_core_030 = ~(input_d[0] | input_c[2]);
  assign cgp_core_031 = input_c[2] ^ input_b[0];
  assign cgp_core_032 = ~(input_a[1] & input_d[0]);
  assign cgp_core_033 = input_b[0] | input_e[1];
  assign cgp_core_034_not = ~input_e[1];
  assign cgp_core_035 = input_e[0] | input_b[2];
  assign cgp_core_037 = ~(input_b[0] & input_c[0]);
  assign cgp_core_038 = input_e[2] & input_b[1];
  assign cgp_core_039 = input_a[2] | input_a[0];
  assign cgp_core_040 = input_a[1] | input_d[0];
  assign cgp_core_042 = input_a[2] & input_b[1];
  assign cgp_core_043 = ~(input_c[0] | input_c[0]);
  assign cgp_core_047 = ~input_e[0];
  assign cgp_core_048 = ~(input_e[0] | input_c[1]);
  assign cgp_core_050 = ~(input_a[1] ^ input_b[1]);
  assign cgp_core_051 = input_d[1] & input_b[0];
  assign cgp_core_055 = input_b[2] | input_e[1];
  assign cgp_core_056 = input_b[1] | input_d[1];
  assign cgp_core_058 = input_a[0] ^ input_c[2];
  assign cgp_core_059 = input_e[2] & input_d[0];
  assign cgp_core_060 = ~(input_a[2] & input_a[0]);
  assign cgp_core_062 = input_a[1] & input_c[0];
  assign cgp_core_064_not = ~input_c[2];
  assign cgp_core_065 = ~(input_c[2] ^ cgp_core_062);
  assign cgp_core_066 = ~input_a[0];
  assign cgp_core_067 = ~(input_e[1] | input_e[0]);
  assign cgp_core_068_not = ~input_d[1];
  assign cgp_core_069 = input_c[1] ^ input_e[0];
  assign cgp_core_070 = input_e[0] & input_d[1];
  assign cgp_core_072 = input_c[0] & input_d[0];
  assign cgp_core_073 = input_d[0] ^ input_d[2];
  assign cgp_core_076 = input_e[1] | input_e[1];
  assign cgp_core_079_not = ~input_c[1];

  assign cgp_out[0] = 1'b0;
endmodule