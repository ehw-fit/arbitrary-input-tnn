module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048_not;
  wire cgp_core_049;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060_not;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_079;

  assign cgp_core_017 = input_g[1] | input_g[0];
  assign cgp_core_019 = input_c[1] ^ input_c[0];
  assign cgp_core_022 = input_d[1] & input_f[1];
  assign cgp_core_023 = ~input_e[0];
  assign cgp_core_024 = ~(input_a[0] ^ input_d[1]);
  assign cgp_core_026 = input_a[1] & input_e[0];
  assign cgp_core_028 = input_b[1] & input_a[1];
  assign cgp_core_030 = input_d[1] | cgp_core_026;
  assign cgp_core_031 = ~(input_f[0] ^ input_c[1]);
  assign cgp_core_032 = ~input_g[0];
  assign cgp_core_034 = input_b[1] | input_c[1];
  assign cgp_core_035 = input_b[1] & input_c[1];
  assign cgp_core_037 = ~(input_e[0] ^ input_f[0]);
  assign cgp_core_039_not = ~input_b[1];
  assign cgp_core_044 = input_g[0] | input_d[0];
  assign cgp_core_045 = ~(input_e[1] ^ input_g[1]);
  assign cgp_core_046 = ~input_g[1];
  assign cgp_core_047 = ~(input_f[0] ^ input_e[1]);
  assign cgp_core_048_not = ~input_a[1];
  assign cgp_core_049 = cgp_core_034 & input_f[1];
  assign cgp_core_050_not = ~input_f[1];
  assign cgp_core_051 = input_g[0] | input_b[1];
  assign cgp_core_053 = ~input_c[1];
  assign cgp_core_055 = input_g[1] | cgp_core_049;
  assign cgp_core_056 = input_g[1] & input_f[1];
  assign cgp_core_057 = cgp_core_035 | cgp_core_056;
  assign cgp_core_058 = ~(input_d[0] & input_g[1]);
  assign cgp_core_060_not = ~cgp_core_057;
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_062 = cgp_core_030 & cgp_core_061;
  assign cgp_core_063 = cgp_core_062 & cgp_core_060_not;
  assign cgp_core_064 = ~(cgp_core_030 ^ cgp_core_055);
  assign cgp_core_065 = cgp_core_064 & cgp_core_060_not;
  assign cgp_core_066 = ~(input_a[1] & input_f[1]);
  assign cgp_core_068 = input_e[1] & cgp_core_065;
  assign cgp_core_069 = ~(input_f[0] ^ input_e[0]);
  assign cgp_core_070 = input_f[1] | input_c[1];
  assign cgp_core_071 = ~(input_g[1] ^ input_b[0]);
  assign cgp_core_074 = ~(input_d[0] | input_g[0]);
  assign cgp_core_079 = cgp_core_068 | cgp_core_063;

  assign cgp_out[0] = cgp_core_079;
endmodule