module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_047_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_070_not;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075_not;
  wire cgp_core_076;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;

  assign cgp_core_018 = input_d[0] ^ input_h[0];
  assign cgp_core_019 = input_g[1] & input_b[0];
  assign cgp_core_021 = input_d[0] & input_a[1];
  assign cgp_core_022 = ~(input_a[0] ^ input_c[0]);
  assign cgp_core_024 = ~(cgp_core_021 ^ input_a[0]);
  assign cgp_core_025 = input_c[0] & cgp_core_018;
  assign cgp_core_026 = ~(input_d[0] & input_h[1]);
  assign cgp_core_028 = input_f[0] | input_f[1];
  assign cgp_core_029 = input_a[0] | input_d[0];
  assign cgp_core_032 = cgp_core_024 ^ input_g[0];
  assign cgp_core_033 = input_b[0] & input_g[0];
  assign cgp_core_034 = input_b[0] ^ input_c[0];
  assign cgp_core_035 = input_a[1] & input_c[0];
  assign cgp_core_036 = input_b[1] ^ input_d[1];
  assign cgp_core_037 = input_b[1] | input_c[1];
  assign cgp_core_038 = cgp_core_036 | input_g[0];
  assign cgp_core_039 = input_a[0] ^ input_h[0];
  assign cgp_core_040 = cgp_core_037 | input_c[1];
  assign cgp_core_043 = ~input_f[1];
  assign cgp_core_044 = input_e[1] & input_g[1];
  assign cgp_core_047_not = ~input_f[0];
  assign cgp_core_049 = input_d[0] & input_h[0];
  assign cgp_core_050 = input_d[0] ^ input_a[1];
  assign cgp_core_052 = input_a[1] ^ input_g[1];
  assign cgp_core_054 = input_g[0] | input_b[0];
  assign cgp_core_055 = input_e[0] ^ cgp_core_054;
  assign cgp_core_057 = input_b[0] ^ input_e[0];
  assign cgp_core_060 = cgp_core_038 & input_f[0];
  assign cgp_core_064 = input_e[0] ^ cgp_core_055;
  assign cgp_core_065 = ~cgp_core_040;
  assign cgp_core_068 = ~cgp_core_065;
  assign cgp_core_069_not = ~input_a[0];
  assign cgp_core_070_not = ~cgp_core_068;
  assign cgp_core_072 = ~input_a[0];
  assign cgp_core_073 = cgp_core_069_not | input_d[0];
  assign cgp_core_075_not = ~input_c[1];
  assign cgp_core_076 = ~(input_d[0] ^ input_b[1]);
  assign cgp_core_079 = input_f[0] & cgp_core_064;
  assign cgp_core_080 = input_d[0] & input_a[1];
  assign cgp_core_081 = input_a[1] ^ cgp_core_064;
  assign cgp_core_083 = ~input_a[1];
  assign cgp_core_084 = input_c[0] & cgp_core_083;
  assign cgp_core_085 = ~(input_g[1] & input_a[0]);
  assign cgp_core_086 = cgp_core_029 ^ input_h[0];
  assign cgp_core_087 = ~input_d[1];
  assign cgp_core_088 = input_b[1] & input_a[1];
  assign cgp_core_089 = ~(cgp_core_025 | input_a[1]);
  assign cgp_core_092 = ~(input_g[1] | cgp_core_087);
  assign cgp_core_093 = ~(cgp_core_085 ^ input_b[1]);
  assign cgp_core_094 = ~input_a[0];

  assign cgp_out[0] = 1'b0;
endmodule