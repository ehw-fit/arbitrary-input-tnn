module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_010;
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041_not;
  wire cgp_core_042;

  assign cgp_core_010 = input_c[0] ^ input_c[0];
  assign cgp_core_011 = input_c[0] & input_d[0];
  assign cgp_core_012 = input_c[1] ^ input_d[1];
  assign cgp_core_013 = input_c[1] | input_d[1];
  assign cgp_core_015 = input_a[1] & input_d[0];
  assign cgp_core_016 = cgp_core_013 | input_a[0];
  assign cgp_core_017 = input_d[1] ^ cgp_core_010;
  assign cgp_core_018 = input_b[0] & cgp_core_010;
  assign cgp_core_019 = input_b[1] | input_d[1];
  assign cgp_core_022 = cgp_core_019 & cgp_core_018;
  assign cgp_core_024 = ~input_d[1];
  assign cgp_core_027 = input_d[0] & input_b[1];
  assign cgp_core_028 = ~(cgp_core_024 & input_a[0]);
  assign cgp_core_030 = ~(input_b[0] | input_a[1]);
  assign cgp_core_031 = cgp_core_018 ^ cgp_core_030;
  assign cgp_core_033 = ~(cgp_core_018 ^ input_a[1]);
  assign cgp_core_034 = ~input_d[0];
  assign cgp_core_036 = cgp_core_017 & input_a[0];
  assign cgp_core_037 = cgp_core_036 & cgp_core_034;
  assign cgp_core_038 = ~(cgp_core_017 ^ input_a[0]);
  assign cgp_core_039 = cgp_core_038 & cgp_core_034;
  assign cgp_core_041_not = ~input_d[1];
  assign cgp_core_042 = ~(cgp_core_027 | cgp_core_041_not);

  assign cgp_out[0] = 1'b1;
endmodule