module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_016_not = ~input_c[1];
  assign cgp_core_017 = input_b[1] ^ input_e[1];
  assign cgp_core_018 = ~(input_a[0] | input_f[1]);
  assign cgp_core_019 = ~(input_b[1] & input_a[0]);
  assign cgp_core_021 = input_b[1] | input_c[1];
  assign cgp_core_022 = input_e[0] & input_a[1];
  assign cgp_core_023 = ~(input_d[0] ^ input_e[1]);
  assign cgp_core_027 = input_b[0] | input_f[1];
  assign cgp_core_028 = ~(input_a[0] & input_c[1]);
  assign cgp_core_031 = input_c[0] & input_f[1];
  assign cgp_core_033 = ~(input_a[1] & input_e[0]);
  assign cgp_core_034 = input_c[1] & input_d[1];
  assign cgp_core_036 = ~input_e[0];
  assign cgp_core_039 = ~(input_f[1] ^ input_e[1]);
  assign cgp_core_040 = ~input_f[1];
  assign cgp_core_041 = input_c[0] & input_b[1];
  assign cgp_core_042 = ~input_e[0];
  assign cgp_core_043 = input_f[1] & input_a[0];
  assign cgp_core_045 = ~(input_e[1] & input_c[1]);
  assign cgp_core_046 = input_d[0] | input_a[1];
  assign cgp_core_047 = input_c[1] | input_a[0];
  assign cgp_core_049 = ~input_f[0];
  assign cgp_core_051 = input_f[1] & input_d[0];
  assign cgp_core_052 = input_f[0] ^ input_e[1];
  assign cgp_core_053 = ~(input_c[1] & input_f[0]);
  assign cgp_core_057 = input_f[1] & input_f[1];
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_061 = ~(input_f[0] & input_c[1]);
  assign cgp_core_064 = input_e[1] ^ input_e[1];
  assign cgp_core_065 = input_a[0] ^ input_a[1];
  assign cgp_core_066 = input_f[1] & input_b[1];
  assign cgp_core_068 = cgp_core_058 | cgp_core_046;
  assign cgp_core_069 = input_d[1] | cgp_core_068;
  assign cgp_core_070 = input_e[1] | input_f[1];
  assign cgp_core_071 = input_c[1] | cgp_core_070;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;

  assign cgp_out[0] = cgp_core_072;
endmodule