module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039_not;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_054;

  assign cgp_core_013 = input_b[1] | input_a[1];
  assign cgp_core_014 = input_b[1] | input_e[1];
  assign cgp_core_015 = input_b[1] & input_a[1];
  assign cgp_core_020 = input_c[0] | input_e[0];
  assign cgp_core_021 = input_a[1] | cgp_core_014;
  assign cgp_core_022 = input_b[0] & input_e[1];
  assign cgp_core_024 = ~(input_e[0] | input_a[0]);
  assign cgp_core_026 = cgp_core_015 | cgp_core_022;
  assign cgp_core_027_not = ~input_d[1];
  assign cgp_core_028 = input_b[1] | input_a[0];
  assign cgp_core_031 = input_c[1] & input_d[1];
  assign cgp_core_035 = input_c[1] ^ input_e[1];
  assign cgp_core_036 = ~(input_d[0] & input_a[0]);
  assign cgp_core_039_not = ~cgp_core_031;
  assign cgp_core_041 = input_e[0] | input_a[0];
  assign cgp_core_043 = cgp_core_021 & cgp_core_039_not;
  assign cgp_core_045 = input_a[1] & input_e[0];
  assign cgp_core_047 = ~(input_c[1] ^ input_a[0]);
  assign cgp_core_048 = ~(input_d[1] | input_e[1]);
  assign cgp_core_050 = input_a[1] ^ input_d[0];
  assign cgp_core_054 = cgp_core_043 | cgp_core_026;

  assign cgp_out[0] = cgp_core_054;
endmodule