module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029_not;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_039;

  assign cgp_core_014 = ~(input_b[1] & input_a[1]);
  assign cgp_core_015 = ~(input_b[1] & input_a[0]);
  assign cgp_core_017 = input_a[2] & input_a[0];
  assign cgp_core_019 = input_a[1] | input_a[0];
  assign cgp_core_020 = input_b[1] & input_c[0];
  assign cgp_core_022_not = ~input_a[1];
  assign cgp_core_023 = ~input_c[0];
  assign cgp_core_024 = ~input_a[2];
  assign cgp_core_025 = ~input_c[2];
  assign cgp_core_026 = input_b[2] & cgp_core_025;
  assign cgp_core_027 = cgp_core_026 & cgp_core_024;
  assign cgp_core_029_not = ~input_b[2];
  assign cgp_core_031 = input_a[0] & input_a[1];
  assign cgp_core_033 = input_a[2] & input_b[2];
  assign cgp_core_035_not = ~input_c[2];
  assign cgp_core_036 = input_b[0] ^ input_a[1];
  assign cgp_core_037_not = ~input_b[1];
  assign cgp_core_039 = input_c[1] ^ input_c[2];

  assign cgp_out[0] = cgp_core_027;
endmodule