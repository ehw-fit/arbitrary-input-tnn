module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_051;
  wire cgp_core_053_not;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = input_f[1] & input_d[0];
  assign cgp_core_019 = ~(input_c[0] ^ input_f[0]);
  assign cgp_core_024 = ~(input_e[0] & input_b[0]);
  assign cgp_core_025 = ~(input_f[0] ^ input_c[1]);
  assign cgp_core_026 = ~(input_e[0] & input_a[1]);
  assign cgp_core_028 = input_b[1] | input_g[1];
  assign cgp_core_030 = ~(input_g[0] | input_g[1]);
  assign cgp_core_031 = input_f[1] | input_f[0];
  assign cgp_core_035 = ~(input_c[1] | input_f[1]);
  assign cgp_core_036 = input_e[1] ^ input_e[0];
  assign cgp_core_037 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_038 = input_b[0] ^ input_b[0];
  assign cgp_core_039 = input_g[0] & input_d[0];
  assign cgp_core_042 = ~(input_b[1] ^ input_d[0]);
  assign cgp_core_043 = ~(input_f[1] ^ input_e[1]);
  assign cgp_core_044 = ~(input_e[0] & input_a[0]);
  assign cgp_core_045 = input_b[0] ^ input_b[0];
  assign cgp_core_046 = input_f[0] ^ input_g[1];
  assign cgp_core_047 = ~input_g[1];
  assign cgp_core_051 = ~(input_d[1] & input_e[1]);
  assign cgp_core_053_not = ~input_g[1];
  assign cgp_core_055 = ~input_c[0];
  assign cgp_core_056 = input_b[0] ^ input_c[0];
  assign cgp_core_057 = ~(input_c[1] | input_f[1]);
  assign cgp_core_058 = input_b[1] ^ input_e[1];
  assign cgp_core_060 = ~(input_b[1] | input_c[1]);
  assign cgp_core_061 = ~(input_b[0] ^ input_g[1]);
  assign cgp_core_062 = ~(input_e[1] & input_g[1]);
  assign cgp_core_063 = input_f[0] | input_b[1];
  assign cgp_core_064 = input_b[0] & input_d[0];
  assign cgp_core_065 = input_d[1] & cgp_core_060;
  assign cgp_core_066 = input_f[0] & input_c[1];
  assign cgp_core_067 = input_d[1] & input_a[0];
  assign cgp_core_068 = input_d[1] ^ input_g[0];
  assign cgp_core_069 = ~input_c[0];
  assign cgp_core_071 = input_e[0] ^ input_f[0];
  assign cgp_core_072 = ~(input_d[1] ^ input_g[1]);
  assign cgp_core_073 = ~(input_e[1] ^ input_g[1]);
  assign cgp_core_074 = ~(input_d[1] & input_c[1]);
  assign cgp_core_075 = input_d[1] ^ input_a[0];
  assign cgp_core_076 = ~(input_g[0] | input_b[0]);
  assign cgp_core_077 = input_c[1] | input_a[1];
  assign cgp_core_078 = ~(input_c[0] ^ input_e[0]);
  assign cgp_core_079 = ~(input_e[0] | input_f[1]);

  assign cgp_out[0] = cgp_core_065;
endmodule