module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_026;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_056_not;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068_not;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_080;

  assign cgp_core_017 = ~input_e[2];
  assign cgp_core_019 = input_a[1] ^ input_a[2];
  assign cgp_core_020 = input_b[1] & input_e[1];
  assign cgp_core_026 = input_b[2] | cgp_core_020;
  assign cgp_core_028_not = ~input_d[2];
  assign cgp_core_029 = input_c[2] & input_c[1];
  assign cgp_core_030 = ~(input_c[2] ^ input_b[1]);
  assign cgp_core_033 = input_d[2] | input_b[1];
  assign cgp_core_034 = input_a[1] & input_d[2];
  assign cgp_core_035_not = ~input_a[2];
  assign cgp_core_036 = input_c[1] | input_e[2];
  assign cgp_core_038 = cgp_core_036 | input_d[2];
  assign cgp_core_040 = ~input_a[0];
  assign cgp_core_041 = input_d[0] | input_d[0];
  assign cgp_core_043 = input_c[1] & input_c[1];
  assign cgp_core_047 = ~(input_e[2] & input_b[1]);
  assign cgp_core_048 = cgp_core_026 | cgp_core_038;
  assign cgp_core_049 = ~(input_a[2] | input_d[0]);
  assign cgp_core_051 = ~(input_c[1] & input_a[2]);
  assign cgp_core_054 = ~input_b[2];
  assign cgp_core_056_not = ~input_e[0];
  assign cgp_core_058 = ~input_e[0];
  assign cgp_core_059 = input_a[1] & input_c[2];
  assign cgp_core_061 = ~input_c[2];
  assign cgp_core_063 = ~cgp_core_048;
  assign cgp_core_064 = input_a[2] & cgp_core_063;
  assign cgp_core_065 = cgp_core_064 & cgp_core_061;
  assign cgp_core_066 = input_d[2] & input_b[2];
  assign cgp_core_068_not = ~input_b[0];
  assign cgp_core_069 = ~(input_d[1] & input_d[0]);
  assign cgp_core_071 = ~(input_c[1] ^ input_d[0]);
  assign cgp_core_072 = input_d[2] & input_e[0];
  assign cgp_core_074 = ~(input_d[1] & input_a[1]);
  assign cgp_core_075 = ~input_c[2];
  assign cgp_core_076 = ~input_c[0];
  assign cgp_core_080 = ~(input_b[2] | input_a[1]);

  assign cgp_out[0] = cgp_core_065;
endmodule