module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060_not;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067_not;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_018 = input_c[1] | input_e[1];
  assign cgp_core_019 = input_c[1] & input_e[1];
  assign cgp_core_021 = cgp_core_018 & input_a[1];
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_023 = ~(input_c[0] & input_g[1]);
  assign cgp_core_024 = ~input_f[1];
  assign cgp_core_026 = input_f[1] | input_b[1];
  assign cgp_core_027 = ~(input_e[1] & input_e[1]);
  assign cgp_core_028 = input_d[0] ^ input_a[1];
  assign cgp_core_029 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_032 = ~input_e[1];
  assign cgp_core_035 = ~(input_b[1] | input_g[1]);
  assign cgp_core_036 = input_d[0] | input_a[1];
  assign cgp_core_037_not = ~input_a[1];
  assign cgp_core_039 = input_d[0] & input_a[1];
  assign cgp_core_041 = input_b[0] & input_a[0];
  assign cgp_core_046 = input_e[1] | input_d[0];
  assign cgp_core_047 = ~input_d[0];
  assign cgp_core_049 = ~(input_c[0] | input_e[1]);
  assign cgp_core_050 = ~input_a[1];
  assign cgp_core_051 = input_c[1] ^ input_e[0];
  assign cgp_core_052 = input_e[0] | input_a[1];
  assign cgp_core_053 = ~(input_g[1] & input_b[0]);
  assign cgp_core_054 = input_b[1] & input_g[1];
  assign cgp_core_055 = ~(input_d[0] ^ input_f[1]);
  assign cgp_core_056 = input_d[1] & input_f[1];
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_060_not = ~cgp_core_057;
  assign cgp_core_062 = input_c[1] & input_g[0];
  assign cgp_core_065 = cgp_core_022 & cgp_core_060_not;
  assign cgp_core_066 = ~(input_e[1] | input_c[0]);
  assign cgp_core_067_not = ~input_c[0];
  assign cgp_core_068 = ~input_e[0];
  assign cgp_core_070 = ~(input_e[1] ^ input_a[1]);
  assign cgp_core_071 = input_a[0] & input_a[1];
  assign cgp_core_072 = ~(input_b[0] ^ input_g[1]);
  assign cgp_core_073 = ~(input_c[1] & input_b[1]);
  assign cgp_core_074 = input_f[1] | input_d[1];
  assign cgp_core_077 = input_c[1] ^ input_a[0];
  assign cgp_core_078 = ~input_b[0];
  assign cgp_core_079 = ~(input_e[1] & input_c[1]);

  assign cgp_out[0] = cgp_core_065;
endmodule