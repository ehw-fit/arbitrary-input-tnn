module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038_not;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056_not;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;

  assign cgp_core_017 = ~(input_c[0] ^ input_b[1]);
  assign cgp_core_018 = input_b[0] | input_a[2];
  assign cgp_core_022 = ~(input_c[0] | input_c[1]);
  assign cgp_core_024 = input_b[2] & input_e[1];
  assign cgp_core_025 = input_d[2] & input_c[1];
  assign cgp_core_027 = ~(input_a[1] | input_a[0]);
  assign cgp_core_031 = input_d[1] ^ input_e[1];
  assign cgp_core_033 = ~(input_e[2] | input_b[1]);
  assign cgp_core_035 = ~(input_b[2] | input_b[1]);
  assign cgp_core_036 = ~(input_c[2] | input_e[2]);
  assign cgp_core_038_not = ~input_b[2];
  assign cgp_core_043 = ~(input_e[0] & input_c[2]);
  assign cgp_core_044 = input_d[2] & input_b[1];
  assign cgp_core_045 = input_b[1] | input_d[1];
  assign cgp_core_049 = ~(input_e[1] & input_d[0]);
  assign cgp_core_051 = ~(input_d[2] & input_a[1]);
  assign cgp_core_054 = input_d[0] ^ input_e[2];
  assign cgp_core_055 = ~(input_c[0] | input_b[1]);
  assign cgp_core_056_not = ~input_b[2];
  assign cgp_core_058 = ~input_e[0];
  assign cgp_core_061 = input_b[2] ^ input_d[0];
  assign cgp_core_062 = ~cgp_core_061;
  assign cgp_core_063 = ~(input_e[1] ^ input_c[1]);
  assign cgp_core_064 = input_a[1] & input_c[1];
  assign cgp_core_065 = input_d[2] ^ input_d[1];
  assign cgp_core_068 = ~cgp_core_045;
  assign cgp_core_069 = ~input_e[2];
  assign cgp_core_071 = ~(input_e[0] & input_b[2]);
  assign cgp_core_072 = input_d[2] | input_e[1];
  assign cgp_core_074 = ~(input_a[0] & input_a[1]);
  assign cgp_core_075 = input_c[0] & input_a[2];
  assign cgp_core_076 = ~(input_b[1] ^ input_d[1]);

  assign cgp_out[0] = 1'b0;
endmodule