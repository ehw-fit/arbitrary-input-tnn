module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058_not;
  wire cgp_core_060_not;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_092;
  wire cgp_core_094;
  wire cgp_core_096;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_020 = input_a[0] | input_d[0];
  assign cgp_core_022 = input_d[0] & input_f[0];
  assign cgp_core_023 = input_a[1] & input_c[1];
  assign cgp_core_025 = ~(input_c[2] | input_b[0]);
  assign cgp_core_026 = cgp_core_023 | input_e[1];
  assign cgp_core_027 = input_c[2] | input_e[2];
  assign cgp_core_028 = input_c[2] & input_e[2];
  assign cgp_core_029 = cgp_core_027 | cgp_core_026;
  assign cgp_core_030 = cgp_core_027 & cgp_core_026;
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = ~input_c[1];
  assign cgp_core_033 = ~input_a[0];
  assign cgp_core_034 = input_e[0] | input_b[1];
  assign cgp_core_035 = input_c[1] & input_e[1];
  assign cgp_core_036 = input_c[2] & input_e[1];
  assign cgp_core_037 = ~input_f[2];
  assign cgp_core_040 = input_a[2] & cgp_core_029;
  assign cgp_core_041 = ~(input_c[2] ^ input_e[2]);
  assign cgp_core_044 = cgp_core_031 | cgp_core_040;
  assign cgp_core_045 = cgp_core_031 & input_a[2];
  assign cgp_core_046 = ~(input_f[0] & input_b[0]);
  assign cgp_core_047 = ~input_b[2];
  assign cgp_core_048 = input_b[2] & input_c[0];
  assign cgp_core_049 = ~input_f[2];
  assign cgp_core_051 = input_e[2] & input_a[1];
  assign cgp_core_052 = ~(input_c[2] & input_e[1]);
  assign cgp_core_053 = ~input_f[0];
  assign cgp_core_054 = input_b[2] & input_f[1];
  assign cgp_core_056 = ~(input_d[2] & input_d[0]);
  assign cgp_core_058_not = ~input_b[2];
  assign cgp_core_060_not = ~input_d[1];
  assign cgp_core_062 = input_a[2] | input_c[2];
  assign cgp_core_064 = input_c[1] ^ input_e[0];
  assign cgp_core_066 = ~(input_a[1] & input_e[2]);
  assign cgp_core_068 = input_f[2] & input_d[2];
  assign cgp_core_070 = cgp_core_054 | cgp_core_068;
  assign cgp_core_074_not = ~input_b[1];
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = cgp_core_044 & cgp_core_075;
  assign cgp_core_078 = input_d[1] | input_e[1];
  assign cgp_core_085 = ~(input_e[2] & input_a[1]);
  assign cgp_core_086 = input_b[2] | input_f[2];
  assign cgp_core_087 = ~(input_d[0] ^ input_a[0]);
  assign cgp_core_089 = ~input_c[2];
  assign cgp_core_092 = input_b[0] | input_f[2];
  assign cgp_core_094 = ~input_b[0];
  assign cgp_core_096 = ~input_a[2];
  assign cgp_core_098 = cgp_core_076 | cgp_core_045;
  assign cgp_core_099 = ~(input_f[2] ^ input_c[1]);

  assign cgp_out[0] = cgp_core_098;
endmodule