module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, input [1:0] input_i, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024_not;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031_not;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_060;
  wire cgp_core_061_not;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071_not;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_088_not;
  wire cgp_core_090_not;
  wire cgp_core_092;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_101;
  wire cgp_core_102;
  wire cgp_core_103;
  wire cgp_core_105;
  wire cgp_core_106;

  assign cgp_core_020 = ~input_h[0];
  assign cgp_core_021 = input_h[0] & input_i[0];
  assign cgp_core_022 = input_b[1] & input_i[1];
  assign cgp_core_023 = input_d[1] & input_i[1];
  assign cgp_core_024_not = ~cgp_core_022;
  assign cgp_core_025 = input_i[1] & input_f[0];
  assign cgp_core_027 = ~(input_a[0] | input_g[0]);
  assign cgp_core_029 = input_d[1] ^ cgp_core_024_not;
  assign cgp_core_030 = input_g[1] & cgp_core_024_not;
  assign cgp_core_031_not = ~cgp_core_029;
  assign cgp_core_036 = input_a[1] ^ input_c[0];
  assign cgp_core_037 = input_h[0] & input_c[0];
  assign cgp_core_038 = input_b[1] | input_c[1];
  assign cgp_core_039 = input_b[1] & input_d[1];
  assign cgp_core_040 = cgp_core_038 ^ cgp_core_037;
  assign cgp_core_041 = input_c[1] & cgp_core_037;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[0] & input_d[1];
  assign cgp_core_045 = input_a[1] ^ input_a[1];
  assign cgp_core_046 = input_a[1] & cgp_core_040;
  assign cgp_core_047 = cgp_core_045 ^ cgp_core_044;
  assign cgp_core_048 = ~(input_f[0] & input_c[0]);
  assign cgp_core_049 = input_i[0] ^ input_h[0];
  assign cgp_core_050 = cgp_core_042 ^ input_f[0];
  assign cgp_core_051 = input_h[0] & input_c[1];
  assign cgp_core_052 = input_f[0] ^ input_b[1];
  assign cgp_core_053 = input_f[0] & input_g[0];
  assign cgp_core_055 = input_f[1] & input_f[0];
  assign cgp_core_060 = ~(input_e[0] | input_b[0]);
  assign cgp_core_061_not = ~input_e[1];
  assign cgp_core_063 = input_d[0] ^ cgp_core_060;
  assign cgp_core_064 = cgp_core_061_not ^ input_h[1];
  assign cgp_core_068 = cgp_core_036 ^ input_a[0];
  assign cgp_core_069 = cgp_core_036 & input_g[1];
  assign cgp_core_071_not = ~input_f[0];
  assign cgp_core_072 = input_i[1] ^ cgp_core_069;
  assign cgp_core_073 = ~(input_e[0] & cgp_core_069);
  assign cgp_core_075 = ~(input_b[1] ^ input_i[0]);
  assign cgp_core_077 = ~(input_g[1] ^ cgp_core_071_not);
  assign cgp_core_078 = input_a[0] & cgp_core_071_not;
  assign cgp_core_088_not = ~input_c[0];
  assign cgp_core_090_not = ~input_i[1];
  assign cgp_core_092 = ~cgp_core_077;
  assign cgp_core_096 = input_e[1] & input_h[1];
  assign cgp_core_097 = cgp_core_072 | input_i[1];
  assign cgp_core_101 = cgp_core_031_not & cgp_core_096;
  assign cgp_core_102 = ~input_g[0];
  assign cgp_core_103 = ~(input_f[1] | cgp_core_102);
  assign cgp_core_105 = ~(cgp_core_027 ^ input_b[1]);
  assign cgp_core_106 = ~(input_i[0] | cgp_core_101);

  assign cgp_out[0] = 1'b0;
endmodule