module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025_not;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074_not;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_099;

  assign cgp_core_021 = input_a[1] & input_d[2];
  assign cgp_core_022 = ~(input_a[1] | input_a[0]);
  assign cgp_core_023 = input_f[0] | input_f[2];
  assign cgp_core_024 = input_a[0] | input_a[0];
  assign cgp_core_025_not = ~input_f[1];
  assign cgp_core_026 = ~input_c[0];
  assign cgp_core_028 = input_f[1] | input_c[2];
  assign cgp_core_030 = ~input_f[0];
  assign cgp_core_031 = input_e[2] | input_c[2];
  assign cgp_core_032 = ~input_a[2];
  assign cgp_core_036 = ~(input_a[2] | input_c[1]);
  assign cgp_core_038 = input_a[1] ^ input_b[1];
  assign cgp_core_039 = ~(input_c[2] & input_a[0]);
  assign cgp_core_040 = input_f[1] & input_f[1];
  assign cgp_core_042 = ~(input_a[0] | input_c[0]);
  assign cgp_core_047 = ~(input_b[0] & input_f[1]);
  assign cgp_core_048 = ~input_b[0];
  assign cgp_core_050 = ~(input_e[1] | input_e[0]);
  assign cgp_core_051 = ~input_e[0];
  assign cgp_core_052 = ~(input_f[1] ^ input_a[0]);
  assign cgp_core_054 = ~(input_f[2] ^ input_b[1]);
  assign cgp_core_056 = ~(input_d[0] | input_d[2]);
  assign cgp_core_057 = ~input_a[2];
  assign cgp_core_058 = ~(input_f[2] ^ input_c[2]);
  assign cgp_core_060 = input_d[2] | input_f[0];
  assign cgp_core_062 = ~(input_e[0] | input_a[1]);
  assign cgp_core_064_not = ~input_c[2];
  assign cgp_core_065 = ~input_d[1];
  assign cgp_core_066 = ~(input_d[2] ^ input_c[1]);
  assign cgp_core_068 = ~(input_e[1] | input_b[2]);
  assign cgp_core_070 = input_a[1] & input_c[1];
  assign cgp_core_071 = input_f[2] & input_b[2];
  assign cgp_core_073 = ~(input_f[2] ^ input_a[2]);
  assign cgp_core_074_not = ~cgp_core_071;
  assign cgp_core_077 = cgp_core_031 & cgp_core_074_not;
  assign cgp_core_078 = ~input_b[1];
  assign cgp_core_080 = input_f[2] | input_d[1];
  assign cgp_core_083 = input_d[2] | input_d[1];
  assign cgp_core_084 = ~input_a[2];
  assign cgp_core_085 = input_e[1] & input_e[0];
  assign cgp_core_086 = input_c[2] & input_a[1];
  assign cgp_core_089 = ~input_a[1];
  assign cgp_core_090 = input_f[0] | input_c[2];
  assign cgp_core_091 = input_e[0] & input_a[1];
  assign cgp_core_092 = input_b[0] ^ input_c[2];
  assign cgp_core_093 = ~input_a[2];
  assign cgp_core_094 = input_c[0] ^ input_f[1];
  assign cgp_core_095 = input_d[0] ^ input_d[0];
  assign cgp_core_096 = ~input_d[2];
  assign cgp_core_097 = ~(input_a[0] ^ input_c[1]);
  assign cgp_core_099 = input_e[0] | input_e[0];

  assign cgp_out[0] = cgp_core_077;
endmodule