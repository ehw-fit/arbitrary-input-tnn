module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_080;

  assign cgp_core_017 = input_d[0] | input_e[0];
  assign cgp_core_018 = input_c[2] | input_a[2];
  assign cgp_core_019 = ~input_d[1];
  assign cgp_core_022 = input_d[1] | input_c[2];
  assign cgp_core_023 = input_a[1] | input_d[1];
  assign cgp_core_024 = ~(input_b[0] | input_c[0]);
  assign cgp_core_028 = input_c[1] & input_e[1];
  assign cgp_core_029_not = ~input_b[2];
  assign cgp_core_030 = ~(input_e[0] | input_d[0]);
  assign cgp_core_033 = ~(input_b[1] | input_d[1]);
  assign cgp_core_034 = input_d[1] & input_a[0];
  assign cgp_core_035 = ~input_e[0];
  assign cgp_core_037 = input_c[2] | input_d[0];
  assign cgp_core_038 = input_a[1] | input_d[1];
  assign cgp_core_039 = ~(input_c[0] ^ input_d[1]);
  assign cgp_core_042 = input_a[2] | input_d[1];
  assign cgp_core_044 = input_c[1] & input_c[1];
  assign cgp_core_045_not = ~input_d[2];
  assign cgp_core_047 = input_b[2] & input_a[2];
  assign cgp_core_049 = input_c[2] & input_a[0];
  assign cgp_core_050 = ~input_c[2];
  assign cgp_core_051 = input_c[1] & input_e[1];
  assign cgp_core_052 = input_b[2] | cgp_core_051;
  assign cgp_core_054 = ~(input_e[0] & input_b[0]);
  assign cgp_core_055 = input_d[2] | cgp_core_052;
  assign cgp_core_057 = input_e[2] | input_c[2];
  assign cgp_core_059 = ~cgp_core_057;
  assign cgp_core_060 = ~(input_a[0] | input_e[0]);
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_062 = cgp_core_061 & cgp_core_059;
  assign cgp_core_064 = ~(input_e[1] | input_e[0]);
  assign cgp_core_065 = ~(input_b[0] | input_e[0]);
  assign cgp_core_067 = input_a[2] & cgp_core_062;
  assign cgp_core_069 = input_e[0] ^ input_b[0];
  assign cgp_core_070 = input_a[1] & cgp_core_067;
  assign cgp_core_071 = ~input_c[0];
  assign cgp_core_072 = cgp_core_071 & cgp_core_067;
  assign cgp_core_073 = input_d[0] ^ input_e[0];
  assign cgp_core_074 = input_a[1] | input_b[1];
  assign cgp_core_075 = ~(input_c[0] ^ input_e[2]);
  assign cgp_core_077 = input_a[0] & cgp_core_072;
  assign cgp_core_080 = cgp_core_070 | cgp_core_077;

  assign cgp_out[0] = cgp_core_080;
endmodule