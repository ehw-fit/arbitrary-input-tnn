module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_093;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;

  assign cgp_core_018 = ~(input_a[1] ^ input_e[0]);
  assign cgp_core_023 = input_g[1] & input_b[1];
  assign cgp_core_024 = input_c[1] | input_b[1];
  assign cgp_core_025 = input_f[0] & input_h[0];
  assign cgp_core_026 = ~(input_e[1] & input_d[0]);
  assign cgp_core_029 = input_c[1] & input_f[1];
  assign cgp_core_030 = input_a[0] ^ input_f[1];
  assign cgp_core_031 = input_d[0] | input_a[1];
  assign cgp_core_032 = cgp_core_024 | cgp_core_031;
  assign cgp_core_033 = cgp_core_024 & cgp_core_031;
  assign cgp_core_034 = input_e[0] | input_a[0];
  assign cgp_core_036 = input_g[1] | input_h[1];
  assign cgp_core_037 = input_g[1] & input_h[1];
  assign cgp_core_041 = ~(input_g[0] & input_h[0]);
  assign cgp_core_042 = ~(input_h[1] & input_d[0]);
  assign cgp_core_043 = input_d[1] | cgp_core_036;
  assign cgp_core_044 = input_d[1] & cgp_core_036;
  assign cgp_core_048 = cgp_core_037 | cgp_core_044;
  assign cgp_core_051 = ~input_d[1];
  assign cgp_core_052 = input_g[0] & input_b[0];
  assign cgp_core_057 = cgp_core_032 | cgp_core_048;
  assign cgp_core_058 = input_a[1] ^ input_c[0];
  assign cgp_core_059 = cgp_core_057 | cgp_core_043;
  assign cgp_core_060 = cgp_core_057 & cgp_core_043;
  assign cgp_core_063 = input_c[1] & input_b[1];
  assign cgp_core_064 = cgp_core_033 | cgp_core_060;
  assign cgp_core_065 = ~(input_g[0] | input_h[0]);
  assign cgp_core_068 = input_b[0] & input_e[1];
  assign cgp_core_069 = ~input_f[0];
  assign cgp_core_070 = input_g[1] & input_b[0];
  assign cgp_core_071 = ~input_h[0];
  assign cgp_core_073 = input_b[0] | input_c[0];
  assign cgp_core_074 = ~input_b[1];
  assign cgp_core_076 = ~(input_e[0] ^ input_g[0]);
  assign cgp_core_078 = ~input_f[1];
  assign cgp_core_079 = cgp_core_059 & cgp_core_078;
  assign cgp_core_081 = ~(cgp_core_059 ^ input_f[1]);
  assign cgp_core_083 = ~input_f[1];
  assign cgp_core_085 = input_a[1] & input_d[0];
  assign cgp_core_086 = ~input_e[1];
  assign cgp_core_087 = cgp_core_086 & cgp_core_081;
  assign cgp_core_088 = input_a[0] | input_c[0];
  assign cgp_core_089 = ~input_h[1];
  assign cgp_core_090 = input_g[0] | input_d[1];
  assign cgp_core_091 = ~(input_d[1] & input_e[1]);
  assign cgp_core_093 = cgp_core_085 | cgp_core_079;
  assign cgp_core_095 = cgp_core_063 | cgp_core_087;
  assign cgp_core_096 = cgp_core_064 | cgp_core_095;
  assign cgp_core_097 = cgp_core_093 | cgp_core_096;

  assign cgp_out[0] = cgp_core_097;
endmodule