module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_098;

  assign cgp_core_020 = input_a[1] ^ input_f[0];
  assign cgp_core_023 = input_a[1] & input_b[1];
  assign cgp_core_024 = input_f[0] ^ input_d[0];
  assign cgp_core_025 = ~(input_d[2] | input_e[0]);
  assign cgp_core_027 = input_a[2] ^ input_b[2];
  assign cgp_core_028 = input_a[2] & input_b[2];
  assign cgp_core_029 = cgp_core_027 ^ cgp_core_023;
  assign cgp_core_030 = cgp_core_027 & cgp_core_023;
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_033 = ~(input_f[1] & input_c[2]);
  assign cgp_core_034 = ~(input_f[0] ^ input_f[1]);
  assign cgp_core_038 = ~(input_a[0] | input_a[0]);
  assign cgp_core_039 = input_c[2] ^ input_d[2];
  assign cgp_core_040 = input_c[2] & input_d[2];
  assign cgp_core_041 = cgp_core_039 ^ input_d[1];
  assign cgp_core_042 = cgp_core_039 & input_d[1];
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;
  assign cgp_core_046 = ~(input_f[0] & input_e[0]);
  assign cgp_core_047 = input_f[1] | input_f[2];
  assign cgp_core_048 = ~input_a[0];
  assign cgp_core_049 = ~(input_f[0] ^ input_f[0]);
  assign cgp_core_050 = input_b[2] & input_a[2];
  assign cgp_core_051 = input_e[2] | input_f[2];
  assign cgp_core_052 = input_e[2] & input_f[2];
  assign cgp_core_053 = cgp_core_051 | input_e[1];
  assign cgp_core_054 = cgp_core_051 & input_e[1];
  assign cgp_core_055 = cgp_core_052 | cgp_core_054;
  assign cgp_core_056 = input_d[2] | input_b[2];
  assign cgp_core_059 = ~(input_e[2] & input_a[0]);
  assign cgp_core_060 = ~(input_b[0] & input_d[1]);
  assign cgp_core_061 = ~(input_e[0] | input_f[1]);
  assign cgp_core_063 = cgp_core_041 ^ cgp_core_053;
  assign cgp_core_064 = cgp_core_041 & cgp_core_053;
  assign cgp_core_065 = cgp_core_063 ^ input_c[1];
  assign cgp_core_066 = cgp_core_063 & input_c[1];
  assign cgp_core_067 = cgp_core_064 | cgp_core_066;
  assign cgp_core_068 = cgp_core_043 | cgp_core_055;
  assign cgp_core_069 = cgp_core_043 & input_e[2];
  assign cgp_core_070 = cgp_core_068 | cgp_core_067;
  assign cgp_core_071 = cgp_core_068 & cgp_core_067;
  assign cgp_core_072 = cgp_core_069 | cgp_core_071;
  assign cgp_core_073 = ~(input_e[0] | input_b[1]);
  assign cgp_core_074 = ~cgp_core_072;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = cgp_core_031 & cgp_core_075;
  assign cgp_core_078 = ~(cgp_core_031 ^ cgp_core_070);
  assign cgp_core_079 = cgp_core_078 & cgp_core_074;
  assign cgp_core_080 = ~cgp_core_065;
  assign cgp_core_081 = cgp_core_029 & cgp_core_080;
  assign cgp_core_082 = cgp_core_081 & cgp_core_079;
  assign cgp_core_083 = ~(cgp_core_029 ^ cgp_core_065);
  assign cgp_core_084 = cgp_core_083 & cgp_core_079;
  assign cgp_core_085 = ~input_f[1];
  assign cgp_core_087 = cgp_core_085 & cgp_core_084;
  assign cgp_core_088 = ~input_d[0];
  assign cgp_core_089 = ~(input_c[1] | input_e[0]);
  assign cgp_core_090 = input_a[2] & input_e[0];
  assign cgp_core_092 = ~(input_d[0] & input_b[2]);
  assign cgp_core_094 = input_d[2] & input_f[2];
  assign cgp_core_095 = cgp_core_087 | cgp_core_082;
  assign cgp_core_098 = cgp_core_095 | cgp_core_076;

  assign cgp_out[0] = cgp_core_098;
endmodule