module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042_not;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060_not;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_016 = ~(input_e[0] ^ input_a[0]);
  assign cgp_core_019 = ~(input_d[1] ^ input_f[1]);
  assign cgp_core_020 = input_a[1] ^ input_d[0];
  assign cgp_core_021 = ~(input_c[1] & input_c[0]);
  assign cgp_core_023 = input_d[0] ^ input_f[0];
  assign cgp_core_024 = ~(input_e[0] | input_e[0]);
  assign cgp_core_025 = input_d[1] | input_g[1];
  assign cgp_core_026 = input_g[1] & input_e[0];
  assign cgp_core_027 = ~(input_c[1] | input_f[0]);
  assign cgp_core_028 = cgp_core_025 & input_c[1];
  assign cgp_core_029 = cgp_core_026 | cgp_core_028;
  assign cgp_core_030 = ~(input_d[0] | input_f[0]);
  assign cgp_core_031 = input_a[1] ^ input_b[1];
  assign cgp_core_032 = input_a[1] & input_c[0];
  assign cgp_core_033_not = ~input_g[1];
  assign cgp_core_034 = input_b[1] ^ input_f[0];
  assign cgp_core_038 = input_d[1] & input_e[1];
  assign cgp_core_040 = input_e[0] ^ input_b[0];
  assign cgp_core_042_not = ~input_c[0];
  assign cgp_core_043 = ~(input_f[1] | input_c[1]);
  assign cgp_core_045 = input_b[1] & input_f[1];
  assign cgp_core_046 = ~(input_g[1] ^ input_g[0]);
  assign cgp_core_051 = ~(input_a[0] | input_d[0]);
  assign cgp_core_052 = input_a[1] & input_b[1];
  assign cgp_core_053 = input_f[1] | input_e[0];
  assign cgp_core_054 = input_f[1] & input_a[1];
  assign cgp_core_055 = cgp_core_052 | cgp_core_054;
  assign cgp_core_056 = cgp_core_045 | cgp_core_055;
  assign cgp_core_057 = cgp_core_045 & input_a[1];
  assign cgp_core_058 = ~input_e[0];
  assign cgp_core_060_not = ~cgp_core_057;
  assign cgp_core_063 = cgp_core_029 & cgp_core_060_not;
  assign cgp_core_064_not = ~cgp_core_056;
  assign cgp_core_068 = input_b[0] | input_a[0];
  assign cgp_core_069 = ~(input_c[1] | input_c[1]);
  assign cgp_core_072 = ~(input_a[1] | input_c[1]);
  assign cgp_core_074 = ~(input_e[1] ^ input_g[1]);
  assign cgp_core_075 = ~(input_e[0] & input_d[1]);
  assign cgp_core_078 = cgp_core_063 | cgp_core_038;
  assign cgp_core_079 = cgp_core_064_not | cgp_core_078;

  assign cgp_out[0] = cgp_core_079;
endmodule