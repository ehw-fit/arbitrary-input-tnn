module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;

  assign cgp_core_014 = ~(input_f[0] ^ input_c[1]);
  assign cgp_core_016 = input_a[1] | input_c[1];
  assign cgp_core_019 = input_d[0] & input_c[0];
  assign cgp_core_020 = input_f[1] | cgp_core_019;
  assign cgp_core_021 = ~(input_a[0] & input_c[0]);
  assign cgp_core_023 = ~input_f[0];
  assign cgp_core_026_not = ~input_b[1];
  assign cgp_core_027 = input_f[1] & input_c[0];
  assign cgp_core_028 = input_c[0] | input_a[1];
  assign cgp_core_029 = input_a[0] ^ input_a[1];
  assign cgp_core_032 = input_e[1] ^ input_d[1];
  assign cgp_core_033 = input_e[0] & input_a[0];
  assign cgp_core_034 = input_d[1] | cgp_core_033;
  assign cgp_core_035 = input_e[1] | cgp_core_034;
  assign cgp_core_036 = input_d[0] & input_d[0];
  assign cgp_core_038 = ~(input_d[1] | input_c[1]);
  assign cgp_core_042 = ~(input_c[1] & input_f[0]);
  assign cgp_core_044 = cgp_core_020 | cgp_core_035;
  assign cgp_core_045 = ~(input_c[1] | input_c[0]);
  assign cgp_core_051 = ~(input_c[0] & input_f[0]);
  assign cgp_core_054 = input_c[1] | input_a[1];
  assign cgp_core_056 = input_d[0] ^ input_f[0];
  assign cgp_core_058 = ~input_c[1];
  assign cgp_core_061 = ~input_b[1];
  assign cgp_core_063 = ~(input_b[1] & input_a[1]);
  assign cgp_core_064 = input_e[1] ^ input_b[1];
  assign cgp_core_067 = input_b[1] ^ input_f[0];
  assign cgp_core_068 = cgp_core_016 | cgp_core_044;
  assign cgp_core_069 = cgp_core_061 | cgp_core_068;
  assign cgp_core_071 = input_c[0] | input_c[1];
  assign cgp_core_072 = ~input_c[1];

  assign cgp_out[0] = cgp_core_069;
endmodule