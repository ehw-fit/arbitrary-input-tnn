module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018_not;
  wire cgp_core_019;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_080;

  assign cgp_core_017 = ~(input_b[2] | input_d[1]);
  assign cgp_core_018_not = ~input_b[2];
  assign cgp_core_019 = input_d[2] | input_e[1];
  assign cgp_core_024 = ~(input_a[2] & input_b[0]);
  assign cgp_core_026 = input_a[1] & input_a[2];
  assign cgp_core_027 = input_e[2] | input_e[0];
  assign cgp_core_029 = ~(input_e[0] ^ input_c[1]);
  assign cgp_core_030 = input_c[2] | input_a[1];
  assign cgp_core_032 = ~input_b[1];
  assign cgp_core_033 = ~input_d[1];
  assign cgp_core_036 = input_d[0] & input_a[0];
  assign cgp_core_037 = ~input_b[2];
  assign cgp_core_038 = ~(input_d[2] | input_e[2]);
  assign cgp_core_039 = ~(input_a[0] ^ input_e[2]);
  assign cgp_core_041 = ~(input_b[1] | input_a[0]);
  assign cgp_core_042 = input_d[1] | input_c[0];
  assign cgp_core_044 = input_a[0] ^ input_b[1];
  assign cgp_core_045 = ~input_a[2];
  assign cgp_core_046 = input_e[2] & input_b[0];
  assign cgp_core_050 = ~input_c[2];
  assign cgp_core_051 = ~input_b[1];
  assign cgp_core_052 = ~(input_c[1] & input_b[1]);
  assign cgp_core_054 = input_b[0] & input_a[0];
  assign cgp_core_055_not = ~input_c[2];
  assign cgp_core_056 = ~(input_b[1] ^ input_c[1]);
  assign cgp_core_057 = ~input_a[0];
  assign cgp_core_059 = ~(input_b[0] & input_b[0]);
  assign cgp_core_060 = ~(input_e[0] & input_a[0]);
  assign cgp_core_063 = input_e[0] & input_e[0];
  assign cgp_core_065 = input_c[2] & input_c[1];
  assign cgp_core_066 = ~(input_a[0] | input_a[0]);
  assign cgp_core_067 = input_a[1] | input_a[2];
  assign cgp_core_068 = ~(input_b[1] | input_c[2]);
  assign cgp_core_070 = ~input_b[1];
  assign cgp_core_072 = ~(input_c[2] ^ input_b[2]);
  assign cgp_core_073 = ~(input_c[1] & input_a[1]);
  assign cgp_core_074 = ~input_b[1];
  assign cgp_core_076 = input_a[2] | input_e[2];
  assign cgp_core_077 = ~input_b[1];
  assign cgp_core_080 = ~(input_b[1] ^ input_c[2]);

  assign cgp_out[0] = cgp_core_038;
endmodule