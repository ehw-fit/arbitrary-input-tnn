module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_033_not;
  wire cgp_core_036_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067_not;
  wire cgp_core_068;
  wire cgp_core_071;
  wire cgp_core_074;

  assign cgp_core_018 = ~(input_a[0] & input_b[0]);
  assign cgp_core_019 = input_a[1] ^ input_c[1];
  assign cgp_core_024 = input_a[2] ^ input_a[2];
  assign cgp_core_025 = ~(input_a[1] | input_c[1]);
  assign cgp_core_026 = cgp_core_024 ^ input_c[1];
  assign cgp_core_028 = ~input_d[0];
  assign cgp_core_033_not = ~input_b[0];
  assign cgp_core_036_not = ~input_b[1];
  assign cgp_core_038 = ~(input_e[0] | input_a[2]);
  assign cgp_core_039 = ~input_b[0];
  assign cgp_core_041 = input_c[2] | input_e[0];
  assign cgp_core_042_not = ~input_c[0];
  assign cgp_core_044 = ~(input_c[0] | cgp_core_033_not);
  assign cgp_core_045 = ~(input_b[0] | input_d[2]);
  assign cgp_core_046 = ~(input_d[2] & input_a[1]);
  assign cgp_core_054 = ~(input_a[0] ^ input_d[2]);
  assign cgp_core_055 = ~input_e[1];
  assign cgp_core_058 = input_c[0] ^ input_a[0];
  assign cgp_core_063 = input_b[2] & input_b[0];
  assign cgp_core_064 = ~cgp_core_063;
  assign cgp_core_065 = ~input_d[2];
  assign cgp_core_066 = ~(cgp_core_065 | input_a[0]);
  assign cgp_core_067_not = ~input_b[0];
  assign cgp_core_068 = ~(input_d[0] & input_e[2]);
  assign cgp_core_071 = input_c[0] & cgp_core_066;
  assign cgp_core_074 = ~input_b[0];

  assign cgp_out[0] = 1'b0;
endmodule