module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_048;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_083_not;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_020 = ~(input_d[0] & input_d[2]);
  assign cgp_core_022_not = ~input_f[2];
  assign cgp_core_023 = input_e[1] & input_a[1];
  assign cgp_core_024 = ~(input_d[1] & input_a[1]);
  assign cgp_core_027 = input_c[2] ^ input_e[2];
  assign cgp_core_028 = input_c[2] & input_e[2];
  assign cgp_core_029 = cgp_core_027 ^ cgp_core_023;
  assign cgp_core_030 = cgp_core_027 & cgp_core_023;
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = ~(input_c[0] & input_c[0]);
  assign cgp_core_035 = ~input_c[0];
  assign cgp_core_038 = ~input_b[0];
  assign cgp_core_039 = input_a[2] ^ cgp_core_029;
  assign cgp_core_040 = input_a[2] & cgp_core_029;
  assign cgp_core_042 = input_e[1] ^ input_a[2];
  assign cgp_core_044 = cgp_core_031 | cgp_core_040;
  assign cgp_core_045 = cgp_core_031 & cgp_core_040;
  assign cgp_core_048 = input_d[0] ^ input_c[0];
  assign cgp_core_052 = input_f[1] | input_b[1];
  assign cgp_core_053 = input_d[2] ^ input_f[2];
  assign cgp_core_054 = input_d[2] & input_f[2];
  assign cgp_core_055 = cgp_core_053 ^ cgp_core_052;
  assign cgp_core_056 = cgp_core_053 & cgp_core_052;
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058 = input_a[2] ^ input_b[1];
  assign cgp_core_059 = ~input_b[0];
  assign cgp_core_060 = input_d[0] & input_a[2];
  assign cgp_core_061 = input_f[1] ^ input_d[2];
  assign cgp_core_065 = input_b[2] ^ cgp_core_055;
  assign cgp_core_066 = input_b[2] & cgp_core_055;
  assign cgp_core_070 = cgp_core_057 | cgp_core_066;
  assign cgp_core_071 = cgp_core_057 & cgp_core_066;
  assign cgp_core_072 = input_a[2] | input_b[1];
  assign cgp_core_074_not = ~cgp_core_071;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = cgp_core_044 & cgp_core_075;
  assign cgp_core_078 = ~(cgp_core_044 ^ cgp_core_070);
  assign cgp_core_079 = cgp_core_078 & cgp_core_074_not;
  assign cgp_core_080 = ~input_d[2];
  assign cgp_core_082 = cgp_core_039 & cgp_core_079;
  assign cgp_core_083_not = ~cgp_core_065;
  assign cgp_core_084 = cgp_core_083_not & cgp_core_079;
  assign cgp_core_085 = ~(input_c[1] | input_c[0]);
  assign cgp_core_088 = ~(input_b[0] & input_e[1]);
  assign cgp_core_090 = input_a[2] ^ input_f[2];
  assign cgp_core_092 = input_d[2] ^ input_e[2];
  assign cgp_core_093 = input_a[2] ^ input_f[2];
  assign cgp_core_094 = input_d[2] ^ input_b[2];
  assign cgp_core_095 = cgp_core_084 | cgp_core_082;
  assign cgp_core_098 = cgp_core_076 | cgp_core_045;
  assign cgp_core_099 = cgp_core_095 | cgp_core_098;

  assign cgp_out[0] = cgp_core_099;
endmodule