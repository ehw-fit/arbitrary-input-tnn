module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016_not;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020_not;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029_not;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_036;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054_not;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;

  assign cgp_core_014 = input_b[0] ^ input_a[1];
  assign cgp_core_015 = ~(input_d[1] & input_b[1]);
  assign cgp_core_016_not = ~input_d[0];
  assign cgp_core_017 = ~(input_c[1] ^ input_e[1]);
  assign cgp_core_018 = input_a[1] | input_d[1];
  assign cgp_core_019 = ~(input_a[0] | input_b[1]);
  assign cgp_core_020_not = ~input_d[0];
  assign cgp_core_023 = input_a[0] | input_a[1];
  assign cgp_core_025 = ~(input_b[1] & input_e[1]);
  assign cgp_core_027 = input_e[1] ^ input_e[0];
  assign cgp_core_028 = input_e[0] ^ input_a[0];
  assign cgp_core_029_not = ~input_f[0];
  assign cgp_core_030 = ~(input_a[0] ^ input_a[0]);
  assign cgp_core_031 = input_b[1] | input_a[1];
  assign cgp_core_036 = ~(input_d[1] & input_e[1]);
  assign cgp_core_040 = input_b[0] & input_f[0];
  assign cgp_core_041 = input_e[1] | cgp_core_040;
  assign cgp_core_042 = input_c[0] ^ input_e[1];
  assign cgp_core_043 = input_d[1] & input_b[1];
  assign cgp_core_044 = input_f[1] | cgp_core_041;
  assign cgp_core_045 = input_f[1] & input_e[1];
  assign cgp_core_046 = cgp_core_043 | cgp_core_045;
  assign cgp_core_048 = ~cgp_core_046;
  assign cgp_core_049 = ~cgp_core_044;
  assign cgp_core_050 = input_a[1] & cgp_core_049;
  assign cgp_core_051 = cgp_core_050 & cgp_core_048;
  assign cgp_core_052 = ~(input_a[1] ^ cgp_core_044);
  assign cgp_core_053 = cgp_core_052 & cgp_core_048;
  assign cgp_core_054_not = ~input_a[1];
  assign cgp_core_055 = input_e[1] | input_c[1];
  assign cgp_core_058 = input_c[0] & cgp_core_053;
  assign cgp_core_059 = input_f[0] & input_a[1];
  assign cgp_core_062 = input_c[1] & input_a[1];
  assign cgp_core_063 = input_c[1] & cgp_core_058;
  assign cgp_core_064 = ~(input_a[0] ^ input_c[0]);
  assign cgp_core_065 = cgp_core_051 | cgp_core_063;
  assign cgp_core_066 = ~(input_b[0] & input_b[0]);

  assign cgp_out[0] = cgp_core_065;
endmodule