module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_055_not;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_080;

  assign cgp_core_017 = ~input_b[0];
  assign cgp_core_018 = ~(input_c[1] & input_d[2]);
  assign cgp_core_020 = ~(input_b[1] | input_c[1]);
  assign cgp_core_021 = input_b[2] & input_c[2];
  assign cgp_core_022 = input_b[0] & input_d[2];
  assign cgp_core_023 = cgp_core_020 ^ input_a[2];
  assign cgp_core_025 = ~(input_b[2] ^ input_e[2]);
  assign cgp_core_026 = input_a[2] | cgp_core_023;
  assign cgp_core_027 = ~(input_a[2] ^ input_b[2]);
  assign cgp_core_030 = input_d[0] & input_e[1];
  assign cgp_core_032 = ~(input_b[0] ^ input_e[1]);
  assign cgp_core_033 = input_a[1] & input_b[2];
  assign cgp_core_034 = input_d[2] ^ input_d[2];
  assign cgp_core_035 = input_d[0] | cgp_core_034;
  assign cgp_core_038 = input_e[2] ^ input_d[1];
  assign cgp_core_041 = ~input_b[2];
  assign cgp_core_049 = cgp_core_026 | cgp_core_038;
  assign cgp_core_051 = ~input_d[2];
  assign cgp_core_055_not = ~input_d[0];
  assign cgp_core_060 = ~cgp_core_055_not;
  assign cgp_core_062 = ~input_b[2];
  assign cgp_core_065 = input_d[2] & input_b[1];
  assign cgp_core_069 = ~(input_b[2] | input_d[0]);
  assign cgp_core_070 = input_b[0] & input_c[2];
  assign cgp_core_073 = ~input_b[1];
  assign cgp_core_076 = ~(input_a[0] & input_d[0]);
  assign cgp_core_078 = input_b[2] & input_b[2];
  assign cgp_core_080 = ~(input_e[1] & input_d[0]);

  assign cgp_out[0] = 1'b0;
endmodule