module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_026_not;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_059_not;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_085;
  wire cgp_core_088;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_096;

  assign cgp_core_021 = input_e[1] & input_b[0];
  assign cgp_core_022 = input_e[1] ^ input_d[1];
  assign cgp_core_023 = ~input_f[0];
  assign cgp_core_026_not = ~cgp_core_023;
  assign cgp_core_027 = ~(input_d[2] | input_a[2]);
  assign cgp_core_029 = ~(input_c[2] & cgp_core_026_not);
  assign cgp_core_030 = input_d[2] & cgp_core_026_not;
  assign cgp_core_032 = input_e[2] | input_d[0];
  assign cgp_core_033 = input_c[0] & input_b[0];
  assign cgp_core_034 = input_c[1] ^ input_d[1];
  assign cgp_core_035 = ~(input_c[1] | input_a[1]);
  assign cgp_core_037 = input_d[2] | input_f[0];
  assign cgp_core_038 = ~(input_e[1] ^ cgp_core_037);
  assign cgp_core_040 = input_c[2] & input_d[1];
  assign cgp_core_044 = input_e[0] ^ input_f[0];
  assign cgp_core_045 = ~(input_e[0] ^ input_f[0]);
  assign cgp_core_046 = input_e[1] ^ input_f[1];
  assign cgp_core_047 = input_e[1] & input_f[1];
  assign cgp_core_049 = cgp_core_046 & cgp_core_045;
  assign cgp_core_050 = input_c[0] | input_f[2];
  assign cgp_core_051 = ~(input_f[0] ^ input_f[2]);
  assign cgp_core_052 = input_f[2] & input_f[2];
  assign cgp_core_053 = cgp_core_051 ^ cgp_core_050;
  assign cgp_core_054 = ~(input_e[2] | cgp_core_050);
  assign cgp_core_055 = ~(input_a[0] ^ cgp_core_054);
  assign cgp_core_056 = cgp_core_032 ^ cgp_core_044;
  assign cgp_core_057 = ~(cgp_core_032 & cgp_core_044);
  assign cgp_core_059_not = ~input_a[1];
  assign cgp_core_060 = input_c[2] ^ cgp_core_057;
  assign cgp_core_061 = input_a[0] | cgp_core_057;
  assign cgp_core_066 = input_d[1] | input_f[0];
  assign cgp_core_067 = input_b[2] | cgp_core_066;
  assign cgp_core_069 = ~(input_c[0] ^ cgp_core_055);
  assign cgp_core_080 = ~input_f[2];
  assign cgp_core_081 = input_f[2] & input_f[1];
  assign cgp_core_082 = input_f[1] & input_b[1];
  assign cgp_core_085 = cgp_core_060 & input_d[0];
  assign cgp_core_088 = ~(input_a[2] | cgp_core_060);
  assign cgp_core_091 = ~(input_a[2] ^ cgp_core_056);
  assign cgp_core_092 = input_e[0] & input_a[2];
  assign cgp_core_096 = cgp_core_092 ^ cgp_core_082;

  assign cgp_out[0] = 1'b0;
endmodule