module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_010;
  wire cgp_core_011;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_027;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041_not;
  wire cgp_core_042;
  wire cgp_core_043;

  assign cgp_core_010 = ~(input_a[0] | input_c[1]);
  assign cgp_core_011 = input_c[1] ^ input_a[0];
  assign cgp_core_014 = ~(input_c[0] & input_b[1]);
  assign cgp_core_015 = ~input_c[0];
  assign cgp_core_016 = input_a[1] & input_d[0];
  assign cgp_core_017 = input_d[1] & input_b[0];
  assign cgp_core_018 = input_d[1] & input_d[1];
  assign cgp_core_019 = ~input_d[0];
  assign cgp_core_021 = ~input_b[0];
  assign cgp_core_024 = ~input_a[1];
  assign cgp_core_027 = input_d[0] ^ input_d[1];
  assign cgp_core_030 = ~input_a[1];
  assign cgp_core_033 = input_b[1] | input_b[1];
  assign cgp_core_035 = ~(input_c[0] ^ input_d[1]);
  assign cgp_core_037 = ~(input_a[0] ^ input_b[1]);
  assign cgp_core_038 = ~(input_a[0] & input_a[1]);
  assign cgp_core_040 = input_c[1] | cgp_core_030;
  assign cgp_core_041_not = ~input_a[1];
  assign cgp_core_042 = input_b[1] | input_d[1];
  assign cgp_core_043 = cgp_core_040 | cgp_core_042;

  assign cgp_out[0] = cgp_core_043;
endmodule