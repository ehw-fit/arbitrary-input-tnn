module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053_not;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_062;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;

  assign cgp_core_016 = input_d[0] ^ input_a[0];
  assign cgp_core_017 = input_d[0] & input_e[0];
  assign cgp_core_018 = ~(input_e[0] ^ input_a[0]);
  assign cgp_core_019 = input_d[1] & input_e[1];
  assign cgp_core_020 = cgp_core_018 ^ input_g[1];
  assign cgp_core_021 = cgp_core_018 & input_c[1];
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_023 = input_a[0] ^ input_a[0];
  assign cgp_core_024 = input_a[0] & cgp_core_016;
  assign cgp_core_025 = input_b[1] ^ cgp_core_020;
  assign cgp_core_026 = input_a[1] & cgp_core_020;
  assign cgp_core_027 = ~(cgp_core_025 & cgp_core_024);
  assign cgp_core_028 = cgp_core_025 | input_c[1];
  assign cgp_core_029 = ~(input_b[1] ^ input_f[0]);
  assign cgp_core_031 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_032 = input_e[1] & input_a[0];
  assign cgp_core_035 = input_b[1] & input_c[0];
  assign cgp_core_038 = input_g[1] | input_a[1];
  assign cgp_core_040 = input_f[0] | input_g[0];
  assign cgp_core_043 = input_b[1] ^ cgp_core_040;
  assign cgp_core_046 = cgp_core_032 ^ input_f[0];
  assign cgp_core_047 = cgp_core_032 | input_f[0];
  assign cgp_core_048 = input_f[0] ^ input_d[0];
  assign cgp_core_049 = input_a[1] & input_f[0];
  assign cgp_core_050 = input_f[1] ^ input_b[0];
  assign cgp_core_053_not = ~cgp_core_038;
  assign cgp_core_054 = ~cgp_core_038;
  assign cgp_core_056 = ~cgp_core_053_not;
  assign cgp_core_057 = ~input_a[1];
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = cgp_core_031 & cgp_core_058;
  assign cgp_core_062 = input_b[0] & input_c[0];
  assign cgp_core_066 = ~cgp_core_050;
  assign cgp_core_067 = input_e[0] & cgp_core_066;
  assign cgp_core_069 = cgp_core_027 & cgp_core_050;
  assign cgp_core_071 = ~cgp_core_046;
  assign cgp_core_074 = ~(cgp_core_023 ^ cgp_core_046);
  assign cgp_core_075 = input_a[1] & input_f[1];
  assign cgp_core_077 = cgp_core_059 | cgp_core_075;

  assign cgp_out[0] = 1'b0;
endmodule