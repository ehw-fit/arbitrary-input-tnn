module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_076;

  assign cgp_core_014 = input_a[10] & input_a[6];
  assign cgp_core_015 = ~input_a[0];
  assign cgp_core_016 = ~(input_a[9] ^ input_a[4]);
  assign cgp_core_017 = ~input_a[6];
  assign cgp_core_020 = input_a[1] | input_a[10];
  assign cgp_core_021 = input_a[0] ^ input_a[4];
  assign cgp_core_022 = ~(input_a[5] ^ input_a[11]);
  assign cgp_core_027 = input_a[7] & input_a[3];
  assign cgp_core_028 = input_a[3] | input_a[4];
  assign cgp_core_031 = input_a[6] & cgp_core_027;
  assign cgp_core_036 = input_a[1] | input_a[1];
  assign cgp_core_038 = ~input_a[2];
  assign cgp_core_040 = ~input_a[11];
  assign cgp_core_041 = input_a[9] & input_a[1];
  assign cgp_core_042 = ~input_a[7];
  assign cgp_core_043 = input_a[0] & cgp_core_041;
  assign cgp_core_044 = ~input_a[6];
  assign cgp_core_049 = input_a[10] & input_a[5];
  assign cgp_core_051 = ~(input_a[7] & input_a[10]);
  assign cgp_core_055 = ~input_a[10];
  assign cgp_core_056 = ~(input_a[6] | input_a[4]);
  assign cgp_core_057 = cgp_core_043 ^ cgp_core_049;
  assign cgp_core_058 = cgp_core_043 & cgp_core_049;
  assign cgp_core_062 = ~(input_a[0] | input_a[7]);
  assign cgp_core_064 = ~(input_a[7] | input_a[8]);
  assign cgp_core_067 = ~(input_a[7] & input_a[1]);
  assign cgp_core_069 = cgp_core_031 ^ cgp_core_057;
  assign cgp_core_070 = cgp_core_031 & cgp_core_057;
  assign cgp_core_071 = ~(input_a[0] | input_a[6]);
  assign cgp_core_076 = cgp_core_058 | cgp_core_070;

  assign cgp_out[0] = input_a[11];
  assign cgp_out[1] = 1'b1;
  assign cgp_out[2] = cgp_core_069;
  assign cgp_out[3] = cgp_core_076;
endmodule