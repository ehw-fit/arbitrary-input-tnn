module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056_not;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_072_not;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;

  assign cgp_core_014 = ~(input_a[8] ^ input_a[4]);
  assign cgp_core_015 = input_a[0] & input_a[6];
  assign cgp_core_016 = ~(input_a[0] & input_a[8]);
  assign cgp_core_017 = input_a[9] ^ input_a[9];
  assign cgp_core_018 = ~(input_a[3] & input_a[7]);
  assign cgp_core_019 = ~(input_a[6] ^ input_a[5]);
  assign cgp_core_023 = ~(input_a[10] & input_a[4]);
  assign cgp_core_024 = input_a[9] & input_a[9];
  assign cgp_core_026 = input_a[1] & input_a[4];
  assign cgp_core_027 = input_a[6] | input_a[3];
  assign cgp_core_029 = input_a[10] ^ input_a[7];
  assign cgp_core_030 = ~(input_a[11] | input_a[1]);
  assign cgp_core_033 = ~(input_a[11] | input_a[9]);
  assign cgp_core_035 = ~(input_a[10] & input_a[2]);
  assign cgp_core_036 = input_a[4] ^ input_a[1];
  assign cgp_core_038 = ~(input_a[9] & input_a[6]);
  assign cgp_core_039 = ~input_a[11];
  assign cgp_core_040 = ~(input_a[6] | input_a[4]);
  assign cgp_core_043 = input_a[4] | input_a[2];
  assign cgp_core_044 = ~(input_a[0] & input_a[6]);
  assign cgp_core_045 = input_a[1] & input_a[10];
  assign cgp_core_046 = input_a[5] ^ input_a[2];
  assign cgp_core_049 = input_a[3] | input_a[2];
  assign cgp_core_051 = ~(input_a[4] & input_a[4]);
  assign cgp_core_052 = ~(input_a[1] | input_a[6]);
  assign cgp_core_054 = input_a[7] ^ input_a[10];
  assign cgp_core_055 = ~input_a[6];
  assign cgp_core_056_not = ~input_a[10];
  assign cgp_core_062 = ~input_a[4];
  assign cgp_core_065 = ~(input_a[2] & input_a[7]);
  assign cgp_core_066 = input_a[9] | input_a[4];
  assign cgp_core_067 = ~(input_a[0] | input_a[3]);
  assign cgp_core_070 = ~(input_a[7] & input_a[10]);
  assign cgp_core_072_not = ~input_a[4];
  assign cgp_core_073 = ~(input_a[2] ^ input_a[8]);
  assign cgp_core_075 = ~(input_a[1] | input_a[1]);
  assign cgp_core_076 = input_a[8] & input_a[7];

  assign cgp_out[0] = input_a[11];
  assign cgp_out[1] = 1'b0;
  assign cgp_out[2] = cgp_core_044;
  assign cgp_out[3] = cgp_core_015;
endmodule