module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_019_not;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_026;
  wire cgp_core_028_not;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034_not;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_040_not;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045_not;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_051;
  wire cgp_core_053_not;

  assign cgp_core_014 = ~(input_e[1] | input_c[1]);
  assign cgp_core_015 = ~input_e[0];
  assign cgp_core_019_not = ~input_c[1];
  assign cgp_core_020 = ~input_a[0];
  assign cgp_core_022 = ~(input_e[1] ^ input_a[1]);
  assign cgp_core_023 = ~input_a[0];
  assign cgp_core_026 = input_c[1] ^ input_c[1];
  assign cgp_core_028_not = ~input_d[0];
  assign cgp_core_030 = input_b[0] ^ input_c[0];
  assign cgp_core_031 = ~(input_b[0] | input_b[1]);
  assign cgp_core_034_not = ~input_b[0];
  assign cgp_core_035 = input_d[0] & input_e[1];
  assign cgp_core_037 = input_c[0] | input_d[1];
  assign cgp_core_040_not = ~input_e[1];
  assign cgp_core_041 = ~input_c[1];
  assign cgp_core_043 = input_d[1] | input_e[1];
  assign cgp_core_044 = ~(input_d[0] ^ input_e[1]);
  assign cgp_core_045_not = ~input_a[0];
  assign cgp_core_046 = ~(input_c[0] & input_c[1]);
  assign cgp_core_047 = ~(input_a[0] ^ cgp_core_026);
  assign cgp_core_048 = ~(input_a[1] | input_c[0]);
  assign cgp_core_051 = input_a[0] | input_e[1];
  assign cgp_core_053_not = ~input_e[1];

  assign cgp_out[0] = 1'b0;
endmodule