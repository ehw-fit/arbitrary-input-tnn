module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, output [0:0] cgp_out);
  wire cgp_core_010;
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_021_not;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;

  assign cgp_core_010 = input_a[0] ^ input_d[0];
  assign cgp_core_011 = ~(input_c[0] | input_c[0]);
  assign cgp_core_012 = ~(input_c[1] & input_c[0]);
  assign cgp_core_013 = input_c[1] & input_d[1];
  assign cgp_core_014 = cgp_core_012 | cgp_core_011;
  assign cgp_core_015 = cgp_core_012 & input_d[0];
  assign cgp_core_016 = cgp_core_013 | input_b[1];
  assign cgp_core_017 = input_b[0] ^ input_b[1];
  assign cgp_core_019 = input_b[1] ^ input_b[0];
  assign cgp_core_021_not = ~input_a[0];
  assign cgp_core_022 = input_b[0] & input_a[1];
  assign cgp_core_024 = cgp_core_016 ^ input_a[1];
  assign cgp_core_028 = cgp_core_024 | input_d[0];
  assign cgp_core_029 = ~cgp_core_028;
  assign cgp_core_030 = ~input_a[0];
  assign cgp_core_031 = cgp_core_021_not & cgp_core_030;
  assign cgp_core_033 = ~input_d[1];
  assign cgp_core_034 = input_d[1] & cgp_core_029;
  assign cgp_core_037 = input_b[0] & input_c[1];
  assign cgp_core_038 = ~cgp_core_017;
  assign cgp_core_039 = ~(cgp_core_038 | input_b[1]);
  assign cgp_core_041 = cgp_core_016 | cgp_core_039;

  assign cgp_out[0] = 1'b1;
endmodule