module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;

  assign cgp_core_014 = input_a[0] ^ input_d[0];
  assign cgp_core_016 = input_d[1] ^ input_c[1];
  assign cgp_core_018 = ~input_c[0];
  assign cgp_core_019 = cgp_core_016 & input_b[1];
  assign cgp_core_021 = input_e[0] ^ input_f[1];
  assign cgp_core_023 = input_e[1] ^ input_f[1];
  assign cgp_core_025 = input_e[0] ^ input_d[1];
  assign cgp_core_026_not = ~cgp_core_023;
  assign cgp_core_028 = input_d[0] ^ cgp_core_021;
  assign cgp_core_029 = input_d[0] & input_f[1];
  assign cgp_core_030 = input_d[1] ^ cgp_core_025;
  assign cgp_core_031 = input_b[1] | cgp_core_025;
  assign cgp_core_032 = input_a[0] ^ cgp_core_029;
  assign cgp_core_038 = ~cgp_core_014;
  assign cgp_core_039 = ~(cgp_core_018 | input_e[1]);
  assign cgp_core_040 = ~(cgp_core_018 | cgp_core_032);
  assign cgp_core_041 = cgp_core_039 ^ cgp_core_038;
  assign cgp_core_042 = input_f[1] ^ input_f[1];
  assign cgp_core_044 = ~(input_f[0] | input_e[1]);
  assign cgp_core_046 = input_e[0] ^ input_f[0];
  assign cgp_core_047 = ~cgp_core_044;
  assign cgp_core_049 = ~(input_b[1] ^ input_f[0]);
  assign cgp_core_050 = ~(input_b[0] ^ input_a[0]);
  assign cgp_core_051 = ~input_f[0];
  assign cgp_core_052 = input_e[0] & cgp_core_051;
  assign cgp_core_053 = ~cgp_core_049;
  assign cgp_core_056 = ~(cgp_core_046 | input_e[1]);
  assign cgp_core_057 = cgp_core_056 ^ input_d[1];
  assign cgp_core_058 = ~input_d[0];
  assign cgp_core_059 = ~(cgp_core_041 ^ cgp_core_058);
  assign cgp_core_060 = cgp_core_059 & cgp_core_057;
  assign cgp_core_061 = ~(input_f[0] ^ input_b[1]);
  assign cgp_core_062 = cgp_core_061 | cgp_core_057;
  assign cgp_core_063 = ~input_b[0];
  assign cgp_core_064 = input_e[1] & cgp_core_063;
  assign cgp_core_066 = ~(input_e[1] ^ input_c[1]);
  assign cgp_core_067 = input_f[1] & cgp_core_062;
  assign cgp_core_068 = ~(input_c[0] | input_c[1]);
  assign cgp_core_070 = input_e[1] | cgp_core_067;
  assign cgp_core_071 = cgp_core_052 | input_f[1];

  assign cgp_out[0] = 1'b1;
endmodule