module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_038_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063_not;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_076;

  assign cgp_core_017 = ~(input_c[2] | input_b[0]);
  assign cgp_core_018 = ~(input_d[2] | input_b[0]);
  assign cgp_core_019 = input_c[2] ^ input_b[1];
  assign cgp_core_020 = input_a[1] & input_b[1];
  assign cgp_core_021 = cgp_core_019 ^ input_b[0];
  assign cgp_core_022 = cgp_core_019 & input_c[0];
  assign cgp_core_023 = input_c[0] | cgp_core_022;
  assign cgp_core_024 = input_a[2] ^ input_b[2];
  assign cgp_core_025 = input_a[2] & input_d[0];
  assign cgp_core_027 = ~(input_e[1] | input_b[0]);
  assign cgp_core_028 = cgp_core_025 | cgp_core_027;
  assign cgp_core_029 = input_d[0] ^ input_b[1];
  assign cgp_core_031 = input_d[1] ^ input_e[1];
  assign cgp_core_032 = ~(input_d[1] | input_b[0]);
  assign cgp_core_033 = ~(input_e[1] & input_e[2]);
  assign cgp_core_038_not = ~input_a[2];
  assign cgp_core_040 = ~input_b[2];
  assign cgp_core_041 = input_e[2] | input_a[2];
  assign cgp_core_042 = input_a[1] & input_e[2];
  assign cgp_core_043 = input_e[1] ^ input_c[2];
  assign cgp_core_044 = input_c[1] & cgp_core_033;
  assign cgp_core_045 = input_d[1] & input_c[1];
  assign cgp_core_046 = cgp_core_043 & cgp_core_042;
  assign cgp_core_047 = input_e[2] | cgp_core_046;
  assign cgp_core_048 = input_b[1] ^ input_a[1];
  assign cgp_core_049 = input_c[2] & input_c[1];
  assign cgp_core_051 = input_c[2] & cgp_core_047;
  assign cgp_core_053 = cgp_core_040 | input_e[0];
  assign cgp_core_054 = cgp_core_040 & input_d[0];
  assign cgp_core_055 = ~cgp_core_054;
  assign cgp_core_056 = ~(cgp_core_054 & input_e[2]);
  assign cgp_core_057 = ~input_a[0];
  assign cgp_core_058 = input_c[0] & cgp_core_057;
  assign cgp_core_061 = input_e[1] ^ cgp_core_056;
  assign cgp_core_062 = cgp_core_048 | input_c[2];
  assign cgp_core_063_not = ~input_d[1];
  assign cgp_core_067 = ~input_c[1];
  assign cgp_core_070 = ~(cgp_core_021 ^ input_d[0]);
  assign cgp_core_071 = input_a[1] & input_d[1];
  assign cgp_core_073 = input_e[2] & input_d[0];
  assign cgp_core_076 = input_c[1] | cgp_core_071;

  assign cgp_out[0] = 1'b0;
endmodule