module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_013;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_050;
  wire cgp_core_054;

  assign cgp_core_013 = ~(input_b[0] | input_a[1]);
  assign cgp_core_015 = input_a[0] ^ input_c[1];
  assign cgp_core_016 = ~input_c[1];
  assign cgp_core_017 = input_d[1] | input_e[1];
  assign cgp_core_019 = ~input_b[1];
  assign cgp_core_021 = ~(input_b[1] ^ input_c[0]);
  assign cgp_core_023 = ~input_a[1];
  assign cgp_core_024 = ~input_c[1];
  assign cgp_core_025 = input_c[1] | input_a[1];
  assign cgp_core_029 = input_a[1] & input_c[1];
  assign cgp_core_031 = input_e[1] | input_e[1];
  assign cgp_core_032 = cgp_core_029 | input_e[1];
  assign cgp_core_034 = cgp_core_025 & cgp_core_032;
  assign cgp_core_035 = input_c[1] | input_a[0];
  assign cgp_core_036 = ~cgp_core_034;
  assign cgp_core_039 = input_d[1] & cgp_core_036;
  assign cgp_core_041 = input_d[0] & cgp_core_036;
  assign cgp_core_044 = input_b[0] & cgp_core_041;
  assign cgp_core_045 = ~(input_d[0] & input_a[0]);
  assign cgp_core_050 = ~(input_e[1] ^ input_c[1]);
  assign cgp_core_054 = cgp_core_044 | cgp_core_039;

  assign cgp_out[0] = cgp_core_054;
endmodule