module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_040;
  wire cgp_core_042_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050_not;
  wire cgp_core_058;
  wire cgp_core_059;

  assign cgp_core_015 = input_c[2] & input_c[1];
  assign cgp_core_017 = input_b[1] ^ input_c[2];
  assign cgp_core_019 = ~input_a[1];
  assign cgp_core_022 = input_a[2] & input_b[2];
  assign cgp_core_023 = ~(input_b[1] ^ input_b[1]);
  assign cgp_core_027 = ~input_d[0];
  assign cgp_core_028 = input_b[1] ^ input_d[2];
  assign cgp_core_029 = input_b[0] | input_d[1];
  assign cgp_core_030 = ~(input_d[0] | input_a[1]);
  assign cgp_core_031 = ~(input_a[1] & input_b[0]);
  assign cgp_core_032 = ~(input_d[1] ^ input_a[0]);
  assign cgp_core_033 = input_a[0] | input_b[1];
  assign cgp_core_034 = ~(input_c[2] & input_a[1]);
  assign cgp_core_035 = ~(input_c[1] & input_d[0]);
  assign cgp_core_036 = ~input_c[2];
  assign cgp_core_040 = ~(input_c[2] | input_d[2]);
  assign cgp_core_042_not = ~input_a[2];
  assign cgp_core_044 = ~(input_c[0] | input_a[0]);
  assign cgp_core_045 = input_b[2] & input_d[1];
  assign cgp_core_047 = input_a[1] ^ input_c[2];
  assign cgp_core_048 = ~(input_d[0] | input_d[0]);
  assign cgp_core_050_not = ~input_a[1];
  assign cgp_core_058 = cgp_core_040 | cgp_core_022;
  assign cgp_core_059 = ~(input_b[2] | input_a[0]);

  assign cgp_out[0] = cgp_core_058;
endmodule