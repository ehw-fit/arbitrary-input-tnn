module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030_not;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_075_not;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_018 = input_b[0] & input_a[0];
  assign cgp_core_019 = ~(input_c[1] & input_b[2]);
  assign cgp_core_021 = ~(cgp_core_019 & input_e[2]);
  assign cgp_core_022 = ~(input_d[0] | cgp_core_018);
  assign cgp_core_023_not = ~cgp_core_022;
  assign cgp_core_024 = ~(input_b[2] & input_d[1]);
  assign cgp_core_025 = ~(input_d[0] & input_e[2]);
  assign cgp_core_028 = input_e[2] | input_c[0];
  assign cgp_core_029 = ~input_d[0];
  assign cgp_core_030_not = ~input_a[0];
  assign cgp_core_033 = input_b[0] | input_c[1];
  assign cgp_core_034 = input_d[1] & cgp_core_030_not;
  assign cgp_core_035 = ~(input_a[1] ^ input_b[1]);
  assign cgp_core_037 = ~(input_b[0] ^ input_a[0]);
  assign cgp_core_039 = ~(input_c[1] & input_e[0]);
  assign cgp_core_040 = input_b[1] | input_b[2];
  assign cgp_core_041 = ~(input_e[2] & cgp_core_029);
  assign cgp_core_042 = input_d[1] & cgp_core_029;
  assign cgp_core_052 = ~input_c[0];
  assign cgp_core_053 = input_b[2] ^ cgp_core_040;
  assign cgp_core_054 = input_e[1] & input_d[2];
  assign cgp_core_056 = cgp_core_053 & cgp_core_052;
  assign cgp_core_057 = ~(input_e[0] ^ cgp_core_056);
  assign cgp_core_058 = ~(input_b[2] & cgp_core_057);
  assign cgp_core_060 = input_d[0] | input_d[0];
  assign cgp_core_061 = ~(input_d[2] & input_a[0]);
  assign cgp_core_062 = input_c[2] & input_e[1];
  assign cgp_core_070 = ~(input_d[2] ^ input_e[0]);
  assign cgp_core_071 = input_d[2] | input_c[0];
  assign cgp_core_075_not = ~input_b[2];
  assign cgp_core_076 = input_e[0] ^ cgp_core_041;
  assign cgp_core_077 = ~input_a[1];
  assign cgp_core_078 = ~cgp_core_070;
  assign cgp_core_079 = input_a[2] | cgp_core_078;
  assign cgp_core_080 = cgp_core_079 | input_a[0];

  assign cgp_out[0] = 1'b0;
endmodule