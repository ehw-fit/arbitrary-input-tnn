module top #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 12,
parameter FEAT_BITS = 3,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1470


)(
    input   [FEAT_CNT * FEAT_BITS   -1:0] features,
    output  [$clog2(CLASS_CNT)      -1:0] prediction
);
localparam  SUM_BITS    = $clog2(HIDDEN_CNT + 1);
localparam  SCORE_BITS  = SUM_BITS + 1;
localparam  INDEX_BITS  = $clog2(FEAT_CNT + 1) + FEAT_BITS;

wire            [FEAT_BITS                  -1:0] feature_array [FEAT_CNT-1:0];
wire            [HIDDEN_CNT                 -1:0] hidden;
wire            [HIDDEN_CNT                 -1:0] hidden_n;
wire            [SUM_BITS                   -1:0] popcount      [CLASS_CNT-1:0]; 
wire            [(SUM_BITS + 1)             -1:0] scores        [CLASS_CNT-1:0]; 
wire            [CLASS_CNT * (SUM_BITS + 1) -1:0] score_vec; 

assign hidden_n = ~hidden;

genvar i;
generate
    for(i=0; i<FEAT_CNT; i=i+1) begin: l1
        assign feature_array[i] = features[i*FEAT_BITS +: FEAT_BITS];
    end
endgenerate
generate
    for(i=0;i<CLASS_CNT;i=i+1) begin: l2
        assign score_vec[i*SCORE_BITS +: SCORE_BITS] = scores[i];
    end
endgenerate



    ltg_0 ltg_0_hn (feature_array[3], feature_array[7], feature_array[10], hidden[0]);
    ltg_1 ltg_1_hn (feature_array[0], feature_array[2], feature_array[6], feature_array[7], feature_array[9], hidden[1]);
    ltg_2 ltg_2_hn (feature_array[0], feature_array[2], hidden[2]);
    ltg_3 ltg_3_hn (feature_array[1], feature_array[2], feature_array[3], feature_array[4], feature_array[9], feature_array[10], hidden[3]);
    ltg_4 ltg_4_hn (feature_array[0], feature_array[1], feature_array[2], feature_array[3], feature_array[8], hidden[4]);
    ltg_5 ltg_5_hn (feature_array[0], feature_array[2], feature_array[4], feature_array[5], feature_array[6], feature_array[9], hidden[5]);
assign hidden[6] = 1;
assign hidden[7] = 0;
    ltg_6 ltg_6_hn (feature_array[3], feature_array[6], feature_array[7], hidden[8]);
    ltg_7 ltg_7_hn (feature_array[2], feature_array[4], feature_array[8], feature_array[9], feature_array[10], hidden[9]);
assign hidden[10] = 0;
    ltg_8 ltg_8_hn (feature_array[1], feature_array[4], feature_array[7], feature_array[10], hidden[11]);
    
    popcount_0 popcount_0_pc ({hidden[11], hidden_n[10], hidden[9], hidden[8], hidden[7], hidden_n[6], hidden[5], hidden[4], hidden[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[0]);
    assign scores[0] = 2*popcount[0] + 0;

    popcount_1 popcount_1_pc ({hidden[11], hidden_n[10], hidden[9], hidden[8], hidden[7], hidden_n[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[1]);
    assign scores[1] = 2*popcount[1] + 0;

    popcount_2 popcount_2_pc ({hidden[11], hidden_n[10], hidden[9], hidden[8], hidden_n[7], hidden[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[2]);
    assign scores[2] = 2*popcount[2] + 0;

    popcount_3 popcount_3_pc ({hidden_n[11], hidden_n[10], hidden[9], hidden[8], hidden_n[7], hidden[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[3]);
    assign scores[3] = 2*popcount[3] + 0;

    popcount_4 popcount_4_pc ({hidden_n[11], hidden_n[10], hidden[9], hidden[8], hidden_n[7], hidden[6], hidden[5], hidden[4], hidden_n[3], hidden_n[2], hidden[1], hidden[0]}, popcount[4]);
    assign scores[4] = 2*popcount[4] + 0;

    popcount_5 popcount_5_pc ({hidden_n[11], hidden[10], hidden[9], hidden_n[8], hidden_n[7], hidden_n[6], hidden[5], hidden_n[4], hidden_n[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[5]);
    assign scores[5] = 2*popcount[5] + 0;

    popcount_6 popcount_6_pc ({hidden_n[11], hidden[10], hidden[9], hidden_n[8], hidden[7], hidden_n[6], hidden[5], hidden[4], hidden[3], hidden_n[2], hidden[1], hidden_n[0]}, popcount[6]);
    assign scores[6] = 2*popcount[6] + 0;



argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS+1)) result (
    .inx(score_vec),
    .outimax(prediction)
);
endmodule
module ltg_0(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, output [0:0] mstc_out);
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_cmp_cmp_gte_i1_3;
  wire mstc_cmp_cmp_gte_pi_3_not;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 = input_0[0] ^ input_2[0];
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0 = input_0[0] & input_2[0];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_0[1] ^ input_2[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 = input_0[1] & input_2[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_0[2] ^ input_2[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 = input_0[2] & input_2[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_cmp_cmp_gte_i1_3 = ~mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  assign mstc_cmp_cmp_gte_pi_3_not = ~mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  assign mstc_cmp_cmp_gte_i1_2 = ~mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_2 = input_1[2] & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_pi_3_not;
  assign mstc_cmp_cmp_gte_pi_2 = ~(input_1[2] ^ mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_pi_3_not;
  assign mstc_cmp_cmp_gte_i1_1 = ~mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_1 = input_1[1] & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(input_1[1] ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_cmp_cmp_gte_and1_0 = input_1[0] & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(input_1[0] ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_and2_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and2_2 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_1(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, input [2:0] input_3, input [2:0] input_4, output [0:0] mstc_out);
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_cmp_cmp_gte_pi_4_not;
  wire mstc_cmp_cmp_gte_i1_3;
  wire mstc_cmp_cmp_gte_and1_3;
  wire mstc_cmp_cmp_gte_and2_3;
  wire mstc_cmp_cmp_gte_pi_3;
  wire mstc_cmp_cmp_gte_psum_3;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 = input_2[0] ^ input_4[0];
  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0 = input_2[0] & input_4[0];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_2[1] ^ input_4[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 = input_2[1] & input_4[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_2[2] ^ input_4[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 = input_2[2] & input_4[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0 = input_1[0] ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0 = input_1[0] & mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0 = input_1[1] ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and0 = input_1[1] & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0 = input_1[2] ^ mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and0 = input_1[2] & mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 = input_0[0] ^ input_3[0];
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0 = input_0[0] & input_3[0];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_0[1] ^ input_3[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 = input_0[1] & input_3[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_0[2] ^ input_3[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 = input_0[2] & input_3[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_cmp_cmp_gte_pi_4_not = ~mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1;
  assign mstc_cmp_cmp_gte_i1_3 = ~mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  assign mstc_cmp_cmp_gte_and1_3 = mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1 & mstc_cmp_cmp_gte_i1_3;
  assign mstc_cmp_cmp_gte_and2_3 = mstc_cmp_cmp_gte_and1_3 & mstc_cmp_cmp_gte_pi_4_not;
  assign mstc_cmp_cmp_gte_pi_3 = ~(mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1 ^ mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0);
  assign mstc_cmp_cmp_gte_psum_3 = mstc_cmp_cmp_gte_pi_3 & mstc_cmp_cmp_gte_pi_4_not;
  assign mstc_cmp_cmp_gte_i1_2 = ~mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_2 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1 & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_pi_2 = ~(mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1 ^ mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_i1_1 = ~mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_1 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1 & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_cmp_cmp_gte_and1_0 = mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0 & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2 = mstc_cmp_cmp_gte_and2_1 | mstc_cmp_cmp_gte_and2_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2 = mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and2_3 | mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_2(input [2:0] input_0, input [2:0] input_1, output [0:0] mstc_out);
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_cmp_cmp_gte_i1_2 = ~input_1[2];
  assign mstc_cmp_cmp_gte_and1_2 = input_0[2] & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_pi_2 = ~(input_0[2] ^ input_1[2]);
  assign mstc_cmp_cmp_gte_i1_1 = ~input_1[1];
  assign mstc_cmp_cmp_gte_and1_1 = input_0[1] & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_pi_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(input_0[1] ^ input_1[1]);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_pi_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~input_1[0];
  assign mstc_cmp_cmp_gte_and1_0 = input_0[0] & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(input_0[0] ^ input_1[0]);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_and2_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and1_2 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_3(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, input [2:0] input_3, input [2:0] input_4, input [2:0] input_5, output [0:0] mstc_out);
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0;
  wire mstc_cmp_cmp_gte_i1_4;
  wire mstc_cmp_cmp_gte_pi_4_not;
  wire mstc_cmp_cmp_gte_i1_3;
  wire mstc_cmp_cmp_gte_and1_3;
  wire mstc_cmp_cmp_gte_and2_3;
  wire mstc_cmp_cmp_gte_pi_3;
  wire mstc_cmp_cmp_gte_psum_3;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 = input_0[0] ^ input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0 = input_0[0] & input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_0[1] ^ input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 = input_0[1] & input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_0[2] ^ input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 = input_0[2] & input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 = input_2[0] ^ input_3[0];
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0 = input_2[0] & input_3[0];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_2[1] ^ input_3[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 = input_2[1] & input_3[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_2[2] ^ input_3[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 = input_2[2] & input_3[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0 = input_4[0] ^ input_5[0];
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0 = input_4[0] & input_5[0];
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 = input_4[1] ^ input_5[1];
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 = input_4[1] & input_5[1];
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 = input_4[2] ^ input_5[2];
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 = input_4[2] & input_5[2];
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0 = mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0 = mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 & mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 & mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 & mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1 = mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0 ^ mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and1 = mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0 & mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0 = mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and0 | mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and1;
  assign mstc_cmp_cmp_gte_i1_4 = ~mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0;
  assign mstc_cmp_cmp_gte_pi_4_not = ~mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0;
  assign mstc_cmp_cmp_gte_i1_3 = ~mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_3 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_cmp_cmp_gte_i1_3;
  assign mstc_cmp_cmp_gte_and2_3 = mstc_cmp_cmp_gte_and1_3 & mstc_cmp_cmp_gte_pi_4_not;
  assign mstc_cmp_cmp_gte_pi_3 = ~(mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_3 = mstc_cmp_cmp_gte_pi_3 & mstc_cmp_cmp_gte_pi_4_not;
  assign mstc_cmp_cmp_gte_i1_2 = ~mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_2 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_pi_2 = ~(mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 ^ mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_i1_1 = ~mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 ^ mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0;
  assign mstc_cmp_cmp_gte_and1_0 = mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 ^ mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2 = mstc_cmp_cmp_gte_and2_1 | mstc_cmp_cmp_gte_and2_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and2_3 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_4(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, input [2:0] input_3, input [2:0] input_4, output [0:0] mstc_out);
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and0;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and1;
  wire mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0;
  wire mstc_cmp_cmp_gte_i1_4;
  wire mstc_cmp_cmp_gte_pi_4_not;
  wire mstc_cmp_cmp_gte_i1_3;
  wire mstc_cmp_cmp_gte_pi_3_not;
  wire mstc_cmp_cmp_gte_psum_3;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 = input_1[0] ^ input_2[0];
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0 = input_1[0] & input_2[0];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_1[1] ^ input_2[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 = input_1[1] & input_2[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_1[2] ^ input_2[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 = input_1[2] & input_2[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0 = input_3[0] ^ input_4[0];
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0 = input_3[0] & input_4[0];
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 = input_3[1] ^ input_4[1];
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 = input_3[1] & input_4[1];
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 = input_3[2] ^ input_4[2];
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 = input_3[2] & input_4[2];
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0 = mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0 = mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 & mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 & mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_3_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_3_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 & mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_3_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_3_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1 = mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0 ^ mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and1 = mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor0 & mstc_neg_sumtree_adder_3_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0 = mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and0 | mstc_neg_sumtree_adder_3_u_rca_fa3_fa_and1;
  assign mstc_cmp_cmp_gte_i1_4 = ~mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0;
  assign mstc_cmp_cmp_gte_pi_4_not = ~mstc_neg_sumtree_adder_3_u_rca_fa3_fa_or0;
  assign mstc_cmp_cmp_gte_i1_3 = ~mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1;
  assign mstc_cmp_cmp_gte_pi_3_not = ~mstc_neg_sumtree_adder_3_u_rca_fa3_fa_xor1;
  assign mstc_cmp_cmp_gte_psum_3 = mstc_cmp_cmp_gte_pi_3_not & mstc_cmp_cmp_gte_pi_4_not;
  assign mstc_cmp_cmp_gte_i1_2 = ~mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_2 = input_0[2] & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_pi_2 = ~(input_0[2] ^ mstc_neg_sumtree_adder_3_u_rca_fa2_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_i1_1 = ~mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_1 = input_0[1] & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(input_0[1] ^ mstc_neg_sumtree_adder_3_u_rca_fa1_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0;
  assign mstc_cmp_cmp_gte_and1_0 = input_0[0] & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(input_0[0] ^ mstc_neg_sumtree_adder_3_u_rca_ha_ha_xor0);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2 = mstc_cmp_cmp_gte_and2_1 | mstc_cmp_cmp_gte_and2_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_psum_0;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_5(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, input [2:0] input_3, input [2:0] input_4, input [2:0] input_5, output [0:0] mstc_out);
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0;
  wire mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1;
  wire mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1;
  wire mstc_cmp_cmp_gte_i1_4;
  wire mstc_cmp_cmp_gte_and1_4;
  wire mstc_cmp_cmp_gte_pi_4;
  wire mstc_cmp_cmp_gte_i1_3;
  wire mstc_cmp_cmp_gte_and1_3;
  wire mstc_cmp_cmp_gte_and2_3;
  wire mstc_cmp_cmp_gte_pi_3;
  wire mstc_cmp_cmp_gte_psum_3;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 = input_2[0] ^ input_4[0];
  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0 = input_2[0] & input_4[0];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_2[1] ^ input_4[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 = input_2[1] & input_4[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_2[2] ^ input_4[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 = input_2[2] & input_4[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0 = input_0[0] ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0 = input_0[0] & mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0 = input_0[1] ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and0 = input_0[1] & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_2_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0 = input_0[2] ^ mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and0 = input_0[2] & mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_2_u_rca_fa2_fa_and1;
  assign mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_pos_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 = input_3[0] ^ input_5[0];
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0 = input_3[0] & input_5[0];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_3[1] ^ input_5[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 = input_3[1] & input_5[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_3[2] ^ input_5[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 = input_3[2] & input_5[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0 = input_1[0] ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0 = input_1[0] & mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 = input_1[1] ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 = input_1[1] & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 = input_1[2] ^ mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 = input_1[2] & mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_cmp_cmp_gte_i1_4 = ~mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1;
  assign mstc_cmp_cmp_gte_and1_4 = mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1 & mstc_cmp_cmp_gte_i1_4;
  assign mstc_cmp_cmp_gte_pi_4 = ~(mstc_pos_sumtree_adder_2_u_rca_fa3_fa_and1 ^ mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1);
  assign mstc_cmp_cmp_gte_i1_3 = ~mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_3 = mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1 & mstc_cmp_cmp_gte_i1_3;
  assign mstc_cmp_cmp_gte_and2_3 = mstc_cmp_cmp_gte_and1_3 & mstc_cmp_cmp_gte_pi_4;
  assign mstc_cmp_cmp_gte_pi_3 = ~(mstc_pos_sumtree_adder_2_u_rca_fa3_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_3 = mstc_cmp_cmp_gte_pi_3 & mstc_cmp_cmp_gte_pi_4;
  assign mstc_cmp_cmp_gte_i1_2 = ~mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_2 = mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1 & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_pi_2 = ~(mstc_pos_sumtree_adder_2_u_rca_fa2_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_i1_1 = ~mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_1 = mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1 & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(mstc_pos_sumtree_adder_2_u_rca_fa1_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  assign mstc_cmp_cmp_gte_and1_0 = mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0 & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(mstc_pos_sumtree_adder_2_u_rca_ha_ha_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2 = mstc_cmp_cmp_gte_and2_1 | mstc_cmp_cmp_gte_and2_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2 = mstc_cmp_cmp_gte_and1_4 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and2_3 | mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_6(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, output [0:0] mstc_out);
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_cmp_cmp_gte_pi_3_not;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 = input_0[0] ^ input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0 = input_0[0] & input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_0[1] ^ input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 = input_0[1] & input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_0[2] ^ input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 = input_0[2] & input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_cmp_cmp_gte_pi_3_not = ~mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0;
  assign mstc_cmp_cmp_gte_i1_2 = ~input_2[2];
  assign mstc_cmp_cmp_gte_and1_2 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_pi_3_not;
  assign mstc_cmp_cmp_gte_pi_2 = ~(mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 ^ input_2[2]);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_pi_3_not;
  assign mstc_cmp_cmp_gte_i1_1 = ~input_2[1];
  assign mstc_cmp_cmp_gte_and1_1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 ^ input_2[1]);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~input_2[0];
  assign mstc_cmp_cmp_gte_and1_0 = mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 ^ input_2[0]);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_and2_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and2_2 | mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_7(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, input [2:0] input_3, input [2:0] input_4, output [0:0] mstc_out);
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1;
  wire mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1;
  wire mstc_cmp_cmp_gte_i1_4;
  wire mstc_cmp_cmp_gte_pi_4_not;
  wire mstc_cmp_cmp_gte_i1_3;
  wire mstc_cmp_cmp_gte_and1_3;
  wire mstc_cmp_cmp_gte_and2_3;
  wire mstc_cmp_cmp_gte_pi_3;
  wire mstc_cmp_cmp_gte_psum_3;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 = input_0[0] ^ input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0 = input_0[0] & input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_0[1] ^ input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 = input_0[1] & input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_0[2] ^ input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 = input_0[2] & input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 = input_3[0] ^ input_4[0];
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0 = input_3[0] & input_4[0];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_3[1] ^ input_4[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 = input_3[1] & input_4[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_3[2] ^ input_4[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 = input_3[2] & input_4[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0 = input_2[0] ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0 = input_2[0] & mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 = input_2[1] ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 = input_2[1] & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 = input_2[2] ^ mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 = input_2[2] & mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_2_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_2_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_neg_sumtree_adder_2_u_rca_fa2_fa_or0;
  assign mstc_cmp_cmp_gte_i1_4 = ~mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1;
  assign mstc_cmp_cmp_gte_pi_4_not = ~mstc_neg_sumtree_adder_2_u_rca_fa3_fa_and1;
  assign mstc_cmp_cmp_gte_i1_3 = ~mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_3 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_cmp_cmp_gte_i1_3;
  assign mstc_cmp_cmp_gte_and2_3 = mstc_cmp_cmp_gte_and1_3 & mstc_cmp_cmp_gte_pi_4_not;
  assign mstc_cmp_cmp_gte_pi_3 = ~(mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_neg_sumtree_adder_2_u_rca_fa3_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_3 = mstc_cmp_cmp_gte_pi_3 & mstc_cmp_cmp_gte_pi_4_not;
  assign mstc_cmp_cmp_gte_i1_2 = ~mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_2 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_pi_2 = ~(mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa2_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_psum_3;
  assign mstc_cmp_cmp_gte_i1_1 = ~mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 ^ mstc_neg_sumtree_adder_2_u_rca_fa1_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0;
  assign mstc_cmp_cmp_gte_and1_0 = mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 ^ mstc_neg_sumtree_adder_2_u_rca_ha_ha_xor0);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2 = mstc_cmp_cmp_gte_and2_1 | mstc_cmp_cmp_gte_and2_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_orred_orreduce_red_XAB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and2_3 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module ltg_8(input [2:0] input_0, input [2:0] input_1, input [2:0] input_2, input [2:0] input_3, output [0:0] mstc_out);
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  wire mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  wire mstc_cmp_cmp_gte_i1_3;
  wire mstc_cmp_cmp_gte_and1_3;
  wire mstc_cmp_cmp_gte_pi_3;
  wire mstc_cmp_cmp_gte_i1_2;
  wire mstc_cmp_cmp_gte_and1_2;
  wire mstc_cmp_cmp_gte_and2_2;
  wire mstc_cmp_cmp_gte_pi_2;
  wire mstc_cmp_cmp_gte_psum_2;
  wire mstc_cmp_cmp_gte_i1_1;
  wire mstc_cmp_cmp_gte_and1_1;
  wire mstc_cmp_cmp_gte_and2_1;
  wire mstc_cmp_cmp_gte_pi_1;
  wire mstc_cmp_cmp_gte_psum_1;
  wire mstc_cmp_cmp_gte_i1_0;
  wire mstc_cmp_cmp_gte_and1_0;
  wire mstc_cmp_cmp_gte_and2_0;
  wire mstc_cmp_cmp_gte_pi_0;
  wire mstc_cmp_cmp_gte_psum_0;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XA_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;
  wire mstc_cmp_cmp_gte_orred_orreduce_red_X_0;

  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 = input_0[0] ^ input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0 = input_0[0] & input_1[0];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_0[1] ^ input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 = input_0[1] & input_1[1];
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_0[2] ^ input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 = input_0[2] & input_1[2];
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_pos_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_pos_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0 = input_2[0] ^ input_3[0];
  assign mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0 = input_2[0] & input_3[0];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 = input_2[1] ^ input_3[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 = input_2[1] & input_3[1];
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_ha_ha_and0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa1_fa_and1;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 = input_2[2] ^ input_3[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 = input_2[2] & input_3[2];
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor0 & mstc_neg_sumtree_adder_1_u_rca_fa1_fa_or0;
  assign mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0 = mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and0 | mstc_neg_sumtree_adder_1_u_rca_fa2_fa_and1;
  assign mstc_cmp_cmp_gte_i1_3 = ~mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0;
  assign mstc_cmp_cmp_gte_and1_3 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 & mstc_cmp_cmp_gte_i1_3;
  assign mstc_cmp_cmp_gte_pi_3 = ~(mstc_pos_sumtree_adder_1_u_rca_fa2_fa_or0 ^ mstc_neg_sumtree_adder_1_u_rca_fa2_fa_or0);
  assign mstc_cmp_cmp_gte_i1_2 = ~mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_2 = mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 & mstc_cmp_cmp_gte_i1_2;
  assign mstc_cmp_cmp_gte_and2_2 = mstc_cmp_cmp_gte_and1_2 & mstc_cmp_cmp_gte_pi_3;
  assign mstc_cmp_cmp_gte_pi_2 = ~(mstc_pos_sumtree_adder_1_u_rca_fa2_fa_xor1 ^ mstc_neg_sumtree_adder_1_u_rca_fa2_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_2 = mstc_cmp_cmp_gte_pi_2 & mstc_cmp_cmp_gte_pi_3;
  assign mstc_cmp_cmp_gte_i1_1 = ~mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1;
  assign mstc_cmp_cmp_gte_and1_1 = mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 & mstc_cmp_cmp_gte_i1_1;
  assign mstc_cmp_cmp_gte_and2_1 = mstc_cmp_cmp_gte_and1_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_pi_1 = ~(mstc_pos_sumtree_adder_1_u_rca_fa1_fa_xor1 ^ mstc_neg_sumtree_adder_1_u_rca_fa1_fa_xor1);
  assign mstc_cmp_cmp_gte_psum_1 = mstc_cmp_cmp_gte_pi_1 & mstc_cmp_cmp_gte_psum_2;
  assign mstc_cmp_cmp_gte_i1_0 = ~mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0;
  assign mstc_cmp_cmp_gte_and1_0 = mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 & mstc_cmp_cmp_gte_i1_0;
  assign mstc_cmp_cmp_gte_and2_0 = mstc_cmp_cmp_gte_and1_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_pi_0 = ~(mstc_pos_sumtree_adder_1_u_rca_ha_ha_xor0 ^ mstc_neg_sumtree_adder_1_u_rca_ha_ha_xor0);
  assign mstc_cmp_cmp_gte_psum_0 = mstc_cmp_cmp_gte_pi_0 & mstc_cmp_cmp_gte_psum_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 = mstc_cmp_cmp_gte_and2_0 | mstc_cmp_cmp_gte_and2_1;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2 = mstc_cmp_cmp_gte_and1_3 | mstc_cmp_cmp_gte_psum_0;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_XB_1 = mstc_cmp_cmp_gte_and2_2 | mstc_cmp_cmp_gte_orred_orreduce_red_XBB_2;
  assign mstc_cmp_cmp_gte_orred_orreduce_red_X_0 = mstc_cmp_cmp_gte_orred_orreduce_red_XA_1 | mstc_cmp_cmp_gte_orred_orreduce_red_XB_1;

  assign mstc_out[0] = mstc_cmp_cmp_gte_orred_orreduce_red_X_0;
endmodule
module popcount_0(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_1(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_2(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_3(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_4(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_5(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module popcount_6(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_014 = input_a[1] ^ input_a[2];
  assign cgp_core_015 = input_a[1] & input_a[2];
  assign cgp_core_016 = input_a[0] ^ cgp_core_014;
  assign cgp_core_017 = input_a[0] & cgp_core_014;
  assign cgp_core_018 = cgp_core_015 | cgp_core_017;
  assign cgp_core_019 = ~input_a[6];
  assign cgp_core_020 = input_a[4] ^ input_a[5];
  assign cgp_core_021 = input_a[4] & input_a[5];
  assign cgp_core_022 = input_a[3] ^ cgp_core_020;
  assign cgp_core_023 = input_a[3] & cgp_core_020;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_026 = cgp_core_016 ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_016 & cgp_core_022;
  assign cgp_core_028 = cgp_core_018 ^ cgp_core_024;
  assign cgp_core_029 = cgp_core_018 & cgp_core_024;
  assign cgp_core_030 = cgp_core_028 ^ cgp_core_027;
  assign cgp_core_031 = cgp_core_028 & cgp_core_027;
  assign cgp_core_032 = cgp_core_029 | cgp_core_031;
  assign cgp_core_034 = ~(input_a[8] & input_a[6]);
  assign cgp_core_036 = ~input_a[5];
  assign cgp_core_038 = input_a[7] ^ input_a[8];
  assign cgp_core_039 = input_a[7] & input_a[8];
  assign cgp_core_040 = input_a[6] ^ cgp_core_038;
  assign cgp_core_041 = input_a[6] & cgp_core_038;
  assign cgp_core_042 = cgp_core_039 | cgp_core_041;
  assign cgp_core_044 = input_a[10] ^ input_a[11];
  assign cgp_core_045 = input_a[10] & input_a[11];
  assign cgp_core_046 = input_a[9] ^ cgp_core_044;
  assign cgp_core_047 = input_a[9] & cgp_core_044;
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_050 = cgp_core_040 ^ cgp_core_046;
  assign cgp_core_051 = cgp_core_040 & cgp_core_046;
  assign cgp_core_052 = cgp_core_042 ^ cgp_core_048;
  assign cgp_core_053 = cgp_core_042 & cgp_core_048;
  assign cgp_core_054 = cgp_core_052 ^ cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_058 = ~(input_a[6] & input_a[4]);
  assign cgp_core_062 = cgp_core_026 ^ cgp_core_050;
  assign cgp_core_063 = cgp_core_026 & cgp_core_050;
  assign cgp_core_064 = cgp_core_030 ^ cgp_core_054;
  assign cgp_core_065 = cgp_core_030 & cgp_core_054;
  assign cgp_core_066 = cgp_core_064 ^ cgp_core_063;
  assign cgp_core_067 = cgp_core_064 & cgp_core_063;
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_069 = cgp_core_032 ^ cgp_core_056;
  assign cgp_core_070 = cgp_core_032 & cgp_core_056;
  assign cgp_core_071 = cgp_core_069 ^ cgp_core_068;
  assign cgp_core_072 = cgp_core_069 & cgp_core_068;
  assign cgp_core_073 = cgp_core_070 | cgp_core_072;
  assign cgp_core_074 = ~input_a[5];
  assign cgp_core_076 = input_a[7] ^ input_a[7];
  assign cgp_core_077 = input_a[1] | input_a[1];
  assign cgp_core_078 = input_a[1] | input_a[6];

  assign cgp_out[0] = cgp_core_062;
  assign cgp_out[1] = cgp_core_066;
  assign cgp_out[2] = cgp_core_071;
  assign cgp_out[3] = cgp_core_073;
endmodule
module argmax #(
    parameter SIZE = 9,
    parameter BITS = 4,
    parameter INDEX_BITS = 4
) (
    input [SIZE*BITS-1:0] inx,
    output [INDEX_BITS-1:0] outimax
);

wire [INDEX_BITS-1:0] interm_argmax [SIZE-1:0];
wire [BITS-1:0] interm_max [SIZE-1:0];

assign interm_max[0] = inx[0+:BITS];
assign interm_argmax[0] = 0;

genvar j;
generate
for (j = 1; j < SIZE; j = j + 1) begin : whatss
	wire huge; //Flag that tracks if current sample is largest so far
	assign huge = inx[j*BITS+:BITS] > interm_max[j-1];
	assign interm_max[j] = huge ? inx[j*BITS+:BITS]:interm_max[j-1]; 
	assign interm_argmax[j] = huge ? j:interm_argmax[j-1];
end
endgenerate

assign outimax = interm_argmax[SIZE-1];

endmodule
