module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_029_not;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;

  assign cgp_core_014 = ~(input_e[0] | input_d[1]);
  assign cgp_core_019 = ~(input_e[1] | input_c[1]);
  assign cgp_core_020 = input_b[0] & input_e[1];
  assign cgp_core_024 = input_b[1] | input_a[0];
  assign cgp_core_025 = ~input_b[0];
  assign cgp_core_026 = input_a[0] | input_d[1];
  assign cgp_core_027 = ~input_c[0];
  assign cgp_core_029_not = ~input_a[1];
  assign cgp_core_031 = ~input_c[0];
  assign cgp_core_032 = input_b[0] | input_c[1];
  assign cgp_core_034 = ~input_a[0];
  assign cgp_core_036 = ~input_c[0];
  assign cgp_core_037 = ~(input_a[0] ^ input_c[1]);
  assign cgp_core_038 = input_c[0] & input_b[0];
  assign cgp_core_041 = input_b[1] & input_c[0];
  assign cgp_core_042 = ~input_b[1];
  assign cgp_core_043 = ~(input_b[0] | input_c[1]);
  assign cgp_core_044 = input_c[1] & input_e[0];
  assign cgp_core_045 = ~input_c[1];
  assign cgp_core_046 = input_e[0] | input_a[0];
  assign cgp_core_047 = input_d[0] ^ input_c[0];
  assign cgp_core_049 = input_d[0] & input_e[0];

  assign cgp_out[0] = 1'b0;
endmodule