module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_078;

  assign cgp_core_016 = input_g[0] ^ input_g[0];
  assign cgp_core_017 = input_e[1] & input_b[1];
  assign cgp_core_018 = input_d[1] | input_e[1];
  assign cgp_core_019 = input_d[1] & input_e[1];
  assign cgp_core_020 = input_e[0] | input_a[0];
  assign cgp_core_021 = cgp_core_018 & input_d[0];
  assign cgp_core_022 = cgp_core_019 | cgp_core_021;
  assign cgp_core_024 = input_d[1] & input_d[0];
  assign cgp_core_026 = input_a[1] & cgp_core_020;
  assign cgp_core_027 = ~(input_d[1] | input_b[0]);
  assign cgp_core_028 = input_e[1] & cgp_core_024;
  assign cgp_core_029 = cgp_core_026 | cgp_core_028;
  assign cgp_core_030 = cgp_core_022 | input_a[1];
  assign cgp_core_031 = cgp_core_022 & cgp_core_029;
  assign cgp_core_032 = ~(input_b[1] & input_g[0]);
  assign cgp_core_033 = ~input_c[1];
  assign cgp_core_034 = input_b[1] | input_c[1];
  assign cgp_core_035 = input_b[1] & input_c[1];
  assign cgp_core_037 = ~(input_e[0] & input_a[0]);
  assign cgp_core_040 = input_g[0] & input_f[0];
  assign cgp_core_041 = input_f[1] | input_g[1];
  assign cgp_core_042 = input_f[1] & input_g[1];
  assign cgp_core_044 = input_c[0] & cgp_core_040;
  assign cgp_core_045 = cgp_core_042 | cgp_core_044;
  assign cgp_core_046 = ~(input_c[0] ^ input_e[1]);
  assign cgp_core_048 = input_a[0] ^ input_a[1];
  assign cgp_core_049 = cgp_core_034 & cgp_core_041;
  assign cgp_core_050 = ~input_c[1];
  assign cgp_core_053 = cgp_core_035 | cgp_core_045;
  assign cgp_core_055 = cgp_core_053 | cgp_core_049;
  assign cgp_core_056 = cgp_core_053 & cgp_core_049;
  assign cgp_core_058 = ~cgp_core_056;
  assign cgp_core_059 = cgp_core_031 & cgp_core_058;
  assign cgp_core_060 = ~input_a[1];
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_062 = cgp_core_030 & cgp_core_061;
  assign cgp_core_065 = input_g[0] | input_d[1];
  assign cgp_core_066 = input_b[0] ^ input_g[0];
  assign cgp_core_069 = ~(input_d[0] | input_c[0]);
  assign cgp_core_070 = ~input_e[0];
  assign cgp_core_071 = input_e[1] ^ input_d[1];
  assign cgp_core_072 = ~(input_f[1] | input_e[0]);
  assign cgp_core_073 = input_f[1] & input_a[1];
  assign cgp_core_074 = ~(input_d[0] & input_a[0]);
  assign cgp_core_076 = input_f[0] & input_f[1];
  assign cgp_core_078 = cgp_core_062 | cgp_core_059;

  assign cgp_out[0] = cgp_core_078;
endmodule