module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019_not;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043_not;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_079;

  assign cgp_core_018 = input_c[1] | input_g[1];
  assign cgp_core_019_not = ~input_c[0];
  assign cgp_core_020 = ~(input_a[1] | input_a[0]);
  assign cgp_core_021 = cgp_core_018 & input_d[0];
  assign cgp_core_023 = input_c[0] & input_g[1];
  assign cgp_core_024 = ~(input_b[0] ^ input_d[1]);
  assign cgp_core_026 = ~(input_a[0] & input_b[0]);
  assign cgp_core_028 = input_d[1] & input_b[0];
  assign cgp_core_029 = ~input_g[0];
  assign cgp_core_030 = ~input_d[0];
  assign cgp_core_032 = input_b[1] | input_d[0];
  assign cgp_core_033 = ~(input_g[1] ^ input_d[1]);
  assign cgp_core_034 = ~(input_f[1] & input_e[1]);
  assign cgp_core_035 = ~(input_e[1] | input_b[1]);
  assign cgp_core_037 = input_c[0] ^ input_a[1];
  assign cgp_core_038 = cgp_core_021 & input_e[0];
  assign cgp_core_039 = ~(input_d[0] ^ input_f[0]);
  assign cgp_core_040 = input_e[1] & input_d[1];
  assign cgp_core_041 = cgp_core_038 | cgp_core_040;
  assign cgp_core_042 = input_c[1] & input_e[1];
  assign cgp_core_043_not = ~input_g[0];
  assign cgp_core_044 = ~(input_e[1] | input_f[0]);
  assign cgp_core_045 = ~(input_b[1] ^ input_c[0]);
  assign cgp_core_046 = ~input_e[1];
  assign cgp_core_048 = ~(input_f[0] ^ input_d[0]);
  assign cgp_core_049 = ~(input_g[0] & input_f[0]);
  assign cgp_core_050 = input_f[1] & input_a[0];
  assign cgp_core_051 = ~(input_e[1] ^ input_c[0]);
  assign cgp_core_053 = ~(input_d[1] ^ input_b[1]);
  assign cgp_core_054 = input_e[0] ^ input_a[0];
  assign cgp_core_055 = ~input_a[0];
  assign cgp_core_056 = ~input_f[0];
  assign cgp_core_058 = ~(input_d[0] ^ input_c[1]);
  assign cgp_core_060 = ~(input_f[1] | input_b[1]);
  assign cgp_core_061 = ~(input_a[1] & input_d[1]);
  assign cgp_core_062 = ~input_g[0];
  assign cgp_core_063 = input_a[1] | input_a[0];
  assign cgp_core_067 = ~(input_f[0] ^ input_e[1]);
  assign cgp_core_069 = input_a[0] ^ input_e[0];
  assign cgp_core_072 = input_c[1] & input_g[1];
  assign cgp_core_075 = ~(input_a[0] | input_f[0]);
  assign cgp_core_076 = cgp_core_072 | cgp_core_060;
  assign cgp_core_079 = cgp_core_076 | cgp_core_041;

  assign cgp_out[0] = cgp_core_079;
endmodule