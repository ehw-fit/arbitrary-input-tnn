module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_030;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045_not;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_059;

  assign cgp_core_015 = input_c[2] | input_b[0];
  assign cgp_core_016 = input_b[1] ^ input_c[1];
  assign cgp_core_019 = input_d[1] ^ input_b[1];
  assign cgp_core_020 = ~(input_b[2] | input_c[2]);
  assign cgp_core_023 = input_c[0] & input_c[2];
  assign cgp_core_024 = input_c[1] ^ input_b[2];
  assign cgp_core_025 = ~(input_a[0] ^ input_c[1]);
  assign cgp_core_026 = input_b[0] & input_b[0];
  assign cgp_core_030 = ~(input_d[1] & input_c[2]);
  assign cgp_core_033 = ~(input_b[1] & input_d[1]);
  assign cgp_core_034 = input_d[2] & input_a[2];
  assign cgp_core_035 = ~input_c[2];
  assign cgp_core_036 = ~(input_a[2] & input_a[2]);
  assign cgp_core_037 = input_d[2] | input_c[2];
  assign cgp_core_038 = ~cgp_core_037;
  assign cgp_core_041 = ~(input_c[1] ^ input_d[1]);
  assign cgp_core_042 = ~(input_a[2] & input_d[2]);
  assign cgp_core_045_not = ~input_d[1];
  assign cgp_core_046 = ~(input_c[2] ^ input_a[0]);
  assign cgp_core_047 = ~(input_a[1] | input_d[2]);
  assign cgp_core_048 = input_d[1] | input_b[0];
  assign cgp_core_050 = ~(input_c[1] ^ input_c[0]);
  assign cgp_core_052 = ~(input_b[0] ^ input_b[0]);
  assign cgp_core_053 = input_a[2] & input_b[2];
  assign cgp_core_059 = cgp_core_053 | cgp_core_038;

  assign cgp_out[0] = cgp_core_059;
endmodule