module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032_not;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_041;

  assign cgp_core_014 = ~(input_c[2] | input_c[1]);
  assign cgp_core_015 = ~(input_a[1] | input_b[2]);
  assign cgp_core_017 = ~(input_a[0] | input_b[1]);
  assign cgp_core_018 = input_a[2] | input_c[2];
  assign cgp_core_019 = input_a[2] & input_c[2];
  assign cgp_core_021 = input_a[0] & input_a[1];
  assign cgp_core_022 = cgp_core_019 | input_c[1];
  assign cgp_core_024 = ~cgp_core_022;
  assign cgp_core_025 = ~cgp_core_018;
  assign cgp_core_026 = input_b[2] & cgp_core_025;
  assign cgp_core_028 = ~(input_c[0] | input_a[1]);
  assign cgp_core_029 = input_b[0] & cgp_core_024;
  assign cgp_core_030 = ~(input_b[0] | input_c[0]);
  assign cgp_core_032_not = ~input_c[2];
  assign cgp_core_034 = input_b[2] & cgp_core_029;
  assign cgp_core_035 = input_a[1] & input_a[0];
  assign cgp_core_036 = ~(input_c[0] & input_c[2]);
  assign cgp_core_038 = ~(input_b[1] ^ input_b[2]);
  assign cgp_core_039 = input_b[1] & cgp_core_034;
  assign cgp_core_041 = cgp_core_026 | cgp_core_039;

  assign cgp_out[0] = cgp_core_041;
endmodule