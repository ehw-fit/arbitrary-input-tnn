module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017_not;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035_not;
  wire cgp_core_036;
  wire cgp_core_037_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_055_not;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074_not;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017_not = ~input_d[0];
  assign cgp_core_018 = input_a[1] | input_e[1];
  assign cgp_core_019 = ~(input_d[0] ^ input_a[0]);
  assign cgp_core_020 = ~input_a[0];
  assign cgp_core_023 = ~input_c[1];
  assign cgp_core_027 = ~(input_a[2] | input_c[0]);
  assign cgp_core_028 = ~input_e[2];
  assign cgp_core_029 = ~(input_a[0] ^ input_a[2]);
  assign cgp_core_030 = ~(input_d[0] ^ input_a[1]);
  assign cgp_core_031 = input_c[1] | input_c[2];
  assign cgp_core_033 = input_d[0] | input_d[2];
  assign cgp_core_035_not = ~input_a[1];
  assign cgp_core_036 = ~(input_c[1] ^ input_e[1]);
  assign cgp_core_037_not = ~input_a[0];
  assign cgp_core_040 = input_b[1] & input_d[1];
  assign cgp_core_041 = input_e[2] | input_b[2];
  assign cgp_core_042 = input_e[2] & input_b[2];
  assign cgp_core_044 = input_d[2] & input_e[0];
  assign cgp_core_045 = input_b[2] & input_e[0];
  assign cgp_core_046 = ~(input_d[1] | input_b[2]);
  assign cgp_core_049 = ~(input_b[2] ^ input_a[2]);
  assign cgp_core_050 = ~input_b[0];
  assign cgp_core_051 = input_a[2] & input_d[2];
  assign cgp_core_055_not = ~input_a[2];
  assign cgp_core_056 = ~cgp_core_051;
  assign cgp_core_057 = cgp_core_041 & cgp_core_056;
  assign cgp_core_061 = input_e[1] ^ input_c[1];
  assign cgp_core_062 = input_e[2] ^ input_d[1];
  assign cgp_core_064 = input_c[1] & input_d[1];
  assign cgp_core_065 = ~input_a[2];
  assign cgp_core_068 = input_d[0] | input_d[0];
  assign cgp_core_069 = input_d[2] & input_b[1];
  assign cgp_core_070 = input_a[0] & input_d[1];
  assign cgp_core_071 = ~(input_d[0] ^ input_d[1]);
  assign cgp_core_074_not = ~input_d[0];
  assign cgp_core_075 = ~(input_b[1] | input_e[0]);
  assign cgp_core_076 = ~(input_b[2] ^ input_d[1]);
  assign cgp_core_077 = input_a[2] | input_a[0];
  assign cgp_core_079 = cgp_core_057 | cgp_core_042;
  assign cgp_core_080 = input_c[2] | cgp_core_079;

  assign cgp_out[0] = cgp_core_080;
endmodule