module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027_not;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072_not;
  wire cgp_core_073;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079_not;
  wire cgp_core_080;

  assign cgp_core_018 = ~(input_d[1] & input_c[0]);
  assign cgp_core_021 = input_a[0] | input_c[2];
  assign cgp_core_024 = ~(input_c[0] | input_d[1]);
  assign cgp_core_026 = ~input_b[2];
  assign cgp_core_027_not = ~input_d[1];
  assign cgp_core_029 = ~(input_c[2] | input_a[0]);
  assign cgp_core_031 = input_d[2] & input_d[1];
  assign cgp_core_032 = ~input_d[2];
  assign cgp_core_035 = input_d[0] ^ input_b[2];
  assign cgp_core_036 = ~(input_c[1] & input_e[1]);
  assign cgp_core_038 = ~(input_d[0] ^ input_d[2]);
  assign cgp_core_042 = input_c[0] ^ input_e[0];
  assign cgp_core_043 = input_c[2] & input_a[2];
  assign cgp_core_048 = input_a[2] ^ input_d[0];
  assign cgp_core_050 = ~(input_e[1] & input_a[0]);
  assign cgp_core_051 = input_a[2] ^ input_a[2];
  assign cgp_core_052 = input_c[1] & input_b[1];
  assign cgp_core_055 = input_c[0] | input_e[0];
  assign cgp_core_056 = input_e[2] ^ input_e[2];
  assign cgp_core_058 = input_a[2] & input_b[2];
  assign cgp_core_059 = cgp_core_058 & input_a[1];
  assign cgp_core_060 = input_b[1] & input_b[0];
  assign cgp_core_061 = input_c[0] | input_c[2];
  assign cgp_core_063 = input_a[1] & input_d[0];
  assign cgp_core_067 = ~(input_b[0] & input_d[2]);
  assign cgp_core_069 = ~(input_c[1] | input_e[0]);
  assign cgp_core_070 = ~(input_a[0] ^ input_a[2]);
  assign cgp_core_072_not = ~input_b[1];
  assign cgp_core_073 = ~(input_c[2] | input_b[0]);
  assign cgp_core_076 = ~(input_d[1] ^ input_c[1]);
  assign cgp_core_078 = input_d[1] ^ input_d[0];
  assign cgp_core_079_not = ~input_e[0];
  assign cgp_core_080 = input_b[2] & input_d[1];

  assign cgp_out[0] = cgp_core_059;
endmodule