module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_081_not;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;

  assign cgp_core_018 = input_b[0] | input_c[0];
  assign cgp_core_019 = input_b[0] & input_c[0];
  assign cgp_core_020 = input_b[1] | input_c[1];
  assign cgp_core_021 = input_b[1] & input_c[1];
  assign cgp_core_023 = cgp_core_020 & cgp_core_019;
  assign cgp_core_024 = cgp_core_021 | cgp_core_023;
  assign cgp_core_025 = input_a[0] ^ cgp_core_018;
  assign cgp_core_026 = input_a[0] & cgp_core_018;
  assign cgp_core_027 = input_c[0] | input_e[1];
  assign cgp_core_028 = ~(input_c[1] & input_c[0]);
  assign cgp_core_029 = input_a[1] | cgp_core_026;
  assign cgp_core_030 = input_a[1] & cgp_core_026;
  assign cgp_core_032 = cgp_core_024 | cgp_core_030;
  assign cgp_core_034 = input_f[1] | input_b[1];
  assign cgp_core_035 = input_g[0] & input_h[0];
  assign cgp_core_036 = input_g[1] | input_h[1];
  assign cgp_core_037 = input_g[1] & input_h[1];
  assign cgp_core_038 = cgp_core_036 | cgp_core_035;
  assign cgp_core_039 = cgp_core_036 & cgp_core_035;
  assign cgp_core_040 = cgp_core_037 | cgp_core_039;
  assign cgp_core_041 = ~(input_f[0] & input_h[1]);
  assign cgp_core_042 = ~(input_a[0] & input_g[0]);
  assign cgp_core_043 = input_d[1] | cgp_core_038;
  assign cgp_core_044 = input_d[1] & cgp_core_038;
  assign cgp_core_048 = cgp_core_040 | cgp_core_044;
  assign cgp_core_049 = input_e[1] & input_a[1];
  assign cgp_core_051 = cgp_core_025 & input_d[0];
  assign cgp_core_052 = cgp_core_029 | cgp_core_043;
  assign cgp_core_053 = cgp_core_029 & cgp_core_043;
  assign cgp_core_054 = cgp_core_052 | cgp_core_051;
  assign cgp_core_055 = cgp_core_052 & cgp_core_051;
  assign cgp_core_056 = cgp_core_053 | cgp_core_055;
  assign cgp_core_057 = cgp_core_032 | cgp_core_048;
  assign cgp_core_058 = input_c[1] ^ input_a[1];
  assign cgp_core_059 = cgp_core_057 | cgp_core_056;
  assign cgp_core_063 = input_b[1] ^ input_d[1];
  assign cgp_core_064 = ~(input_h[1] ^ input_g[1]);
  assign cgp_core_065 = ~(input_c[1] & input_b[0]);
  assign cgp_core_067 = ~input_d[0];
  assign cgp_core_070 = input_e[1] & input_f[1];
  assign cgp_core_071 = ~(input_f[1] | input_h[0]);
  assign cgp_core_072 = ~(input_f[1] & input_d[1]);
  assign cgp_core_075 = ~(input_d[0] & input_g[1]);
  assign cgp_core_077 = input_c[0] & input_g[0];
  assign cgp_core_081_not = ~cgp_core_070;
  assign cgp_core_083 = ~input_f[0];
  assign cgp_core_085 = cgp_core_054 & cgp_core_081_not;
  assign cgp_core_086 = ~(input_e[1] | input_f[1]);
  assign cgp_core_088 = input_g[0] & input_g[0];
  assign cgp_core_089 = ~(input_d[1] | input_h[0]);
  assign cgp_core_091 = ~input_b[0];
  assign cgp_core_092 = input_d[1] | input_h[0];
  assign cgp_core_093 = cgp_core_085 | cgp_core_059;
  assign cgp_core_094 = cgp_core_086 | cgp_core_093;
  assign cgp_core_095 = ~(input_h[1] ^ input_g[1]);
  assign cgp_core_096 = input_h[0] | input_c[1];
  assign cgp_core_097 = ~(input_c[0] ^ input_f[1]);

  assign cgp_out[0] = cgp_core_094;
endmodule