module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060_not;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_g[1] & input_e[0]);
  assign cgp_core_018 = input_c[1] | input_e[1];
  assign cgp_core_019 = input_c[1] & input_e[1];
  assign cgp_core_021 = ~input_d[0];
  assign cgp_core_023 = input_d[0] | input_c[1];
  assign cgp_core_025 = input_d[0] | input_e[1];
  assign cgp_core_026 = input_a[1] & cgp_core_018;
  assign cgp_core_027 = input_c[1] | input_e[0];
  assign cgp_core_028 = input_a[0] ^ input_b[0];
  assign cgp_core_030 = cgp_core_019 | cgp_core_026;
  assign cgp_core_031 = ~(input_e[1] | input_f[0]);
  assign cgp_core_033 = input_g[1] & input_e[0];
  assign cgp_core_035 = input_d[1] & input_f[0];
  assign cgp_core_036 = ~(input_f[0] | input_a[1]);
  assign cgp_core_038 = cgp_core_035 | input_g[1];
  assign cgp_core_040 = input_a[1] | input_b[0];
  assign cgp_core_041 = input_b[0] | input_g[0];
  assign cgp_core_042 = input_f[1] & input_b[1];
  assign cgp_core_046 = input_f[0] ^ input_f[0];
  assign cgp_core_048 = ~(input_b[0] | input_d[0]);
  assign cgp_core_049 = input_b[1] | input_f[0];
  assign cgp_core_052 = input_b[1] | input_f[1];
  assign cgp_core_053 = cgp_core_038 | cgp_core_042;
  assign cgp_core_054 = ~(input_f[0] | input_d[0]);
  assign cgp_core_055 = input_d[0] | input_d[1];
  assign cgp_core_056 = cgp_core_053 & cgp_core_052;
  assign cgp_core_058 = input_b[1] ^ input_f[0];
  assign cgp_core_059 = input_b[1] ^ input_g[0];
  assign cgp_core_060_not = ~cgp_core_056;
  assign cgp_core_063 = cgp_core_030 & cgp_core_060_not;
  assign cgp_core_064 = ~(input_f[1] | cgp_core_055);
  assign cgp_core_066 = input_b[0] & input_a[1];
  assign cgp_core_068 = input_a[1] & cgp_core_064;
  assign cgp_core_070 = ~input_a[0];
  assign cgp_core_072 = input_d[1] ^ input_c[1];
  assign cgp_core_073 = input_d[0] & input_a[1];
  assign cgp_core_074 = input_c[0] | input_a[1];
  assign cgp_core_077 = input_f[1] ^ input_c[1];
  assign cgp_core_079 = cgp_core_068 | cgp_core_063;

  assign cgp_out[0] = cgp_core_079;
endmodule