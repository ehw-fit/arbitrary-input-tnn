module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_058;
  wire cgp_core_059_not;

  assign cgp_core_018 = ~(input_a[1] | input_d[1]);
  assign cgp_core_019 = ~(input_c[0] & input_a[1]);
  assign cgp_core_020 = input_c[0] | input_c[2];
  assign cgp_core_022 = ~(input_b[1] | input_b[2]);
  assign cgp_core_025 = ~(input_b[0] | input_b[0]);
  assign cgp_core_026 = input_a[2] ^ input_a[2];
  assign cgp_core_027 = ~(input_d[0] ^ input_d[0]);
  assign cgp_core_028 = ~(input_a[2] ^ input_b[0]);
  assign cgp_core_029 = input_d[0] & input_c[1];
  assign cgp_core_030 = ~(input_d[2] ^ input_d[0]);
  assign cgp_core_031 = input_d[1] | input_d[1];
  assign cgp_core_033 = ~input_d[1];
  assign cgp_core_034 = input_b[1] ^ input_d[0];
  assign cgp_core_036 = ~(input_b[2] ^ input_d[2]);
  assign cgp_core_038 = ~input_d[2];
  assign cgp_core_039 = input_b[2] & cgp_core_038;
  assign cgp_core_042 = ~(input_d[0] | input_d[0]);
  assign cgp_core_047 = input_d[1] & input_c[1];
  assign cgp_core_049 = ~(input_b[1] | input_c[1]);
  assign cgp_core_052 = input_c[2] ^ input_b[2];
  assign cgp_core_053 = ~(input_b[2] & input_b[2]);
  assign cgp_core_054 = ~(input_c[2] ^ input_d[0]);
  assign cgp_core_055 = input_c[1] ^ input_a[1];
  assign cgp_core_058 = input_a[2] | cgp_core_039;
  assign cgp_core_059_not = ~input_c[1];

  assign cgp_out[0] = cgp_core_058;
endmodule