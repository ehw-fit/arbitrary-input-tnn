module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_044_not;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057_not;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063_not;
  wire cgp_core_065;

  assign cgp_core_016 = input_a[1] ^ input_c[1];
  assign cgp_core_019 = ~(cgp_core_016 | input_a[0]);
  assign cgp_core_021 = input_b[0] ^ input_d[0];
  assign cgp_core_023 = input_c[0] ^ input_d[0];
  assign cgp_core_024 = input_b[1] | input_d[1];
  assign cgp_core_025 = cgp_core_023 ^ input_a[0];
  assign cgp_core_026 = cgp_core_023 & input_a[1];
  assign cgp_core_027 = ~(cgp_core_024 & cgp_core_026);
  assign cgp_core_028 = ~(input_e[0] | input_f[0]);
  assign cgp_core_029 = input_e[0] & input_f[0];
  assign cgp_core_031 = input_a[0] & input_e[0];
  assign cgp_core_032 = ~(input_c[0] & cgp_core_029);
  assign cgp_core_034 = ~(input_f[1] ^ input_c[1]);
  assign cgp_core_035 = input_d[1] ^ cgp_core_028;
  assign cgp_core_036 = input_a[0] & input_d[1];
  assign cgp_core_037 = ~input_d[0];
  assign cgp_core_038 = cgp_core_025 | input_e[1];
  assign cgp_core_039 = cgp_core_037 ^ input_c[0];
  assign cgp_core_040 = input_e[1] & input_b[0];
  assign cgp_core_042 = cgp_core_027 ^ input_b[0];
  assign cgp_core_044_not = ~input_f[1];
  assign cgp_core_045 = ~cgp_core_042;
  assign cgp_core_046 = input_b[1] | input_e[1];
  assign cgp_core_047 = input_d[1] & input_c[1];
  assign cgp_core_048 = ~cgp_core_046;
  assign cgp_core_049 = ~input_b[0];
  assign cgp_core_050 = input_a[1] & input_b[1];
  assign cgp_core_051 = cgp_core_050 & cgp_core_048;
  assign cgp_core_053 = ~input_a[0];
  assign cgp_core_054 = ~(input_e[0] & input_c[1]);
  assign cgp_core_055 = input_d[0] & input_c[0];
  assign cgp_core_056 = input_e[1] & input_f[0];
  assign cgp_core_057_not = ~cgp_core_039;
  assign cgp_core_059 = ~cgp_core_035;
  assign cgp_core_060 = input_a[0] & input_b[0];
  assign cgp_core_063_not = ~input_d[1];
  assign cgp_core_065 = cgp_core_051 | input_d[1];

  assign cgp_out[0] = input_c[1];
endmodule