module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_025_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_036_not;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;

  assign cgp_core_017 = input_d[0] & input_e[0];
  assign cgp_core_018 = input_d[1] & input_e[1];
  assign cgp_core_019 = input_d[1] & input_e[1];
  assign cgp_core_021 = ~cgp_core_018;
  assign cgp_core_022 = cgp_core_019 | input_e[0];
  assign cgp_core_023 = input_a[0] ^ input_f[1];
  assign cgp_core_025_not = ~input_a[1];
  assign cgp_core_028 = cgp_core_025_not & input_a[0];
  assign cgp_core_029 = ~(input_a[0] | input_a[0]);
  assign cgp_core_030 = ~cgp_core_022;
  assign cgp_core_031 = cgp_core_022 & input_e[1];
  assign cgp_core_034 = input_b[1] ^ input_f[1];
  assign cgp_core_035 = input_b[1] & input_f[0];
  assign cgp_core_036_not = ~cgp_core_034;
  assign cgp_core_038 = cgp_core_035 | cgp_core_034;
  assign cgp_core_039 = input_f[0] ^ input_g[0];
  assign cgp_core_040 = input_f[0] & input_g[0];
  assign cgp_core_042 = input_b[0] | input_g[1];
  assign cgp_core_046 = ~(input_c[1] ^ cgp_core_039);
  assign cgp_core_048 = input_c[0] ^ input_c[1];
  assign cgp_core_049 = input_c[1] & input_e[0];
  assign cgp_core_050 = input_d[0] ^ input_g[0];
  assign cgp_core_052 = cgp_core_049 | input_a[0];
  assign cgp_core_054 = ~(cgp_core_038 & cgp_core_042);
  assign cgp_core_055 = input_e[0] ^ cgp_core_052;
  assign cgp_core_057 = input_f[0] | input_g[0];
  assign cgp_core_058 = ~cgp_core_057;
  assign cgp_core_059 = input_e[1] & cgp_core_058;
  assign cgp_core_061 = ~(cgp_core_055 ^ cgp_core_055);
  assign cgp_core_062 = input_e[1] & input_f[0];
  assign cgp_core_063 = ~cgp_core_062;
  assign cgp_core_066 = ~input_d[0];
  assign cgp_core_067 = ~input_a[0];
  assign cgp_core_069_not = ~cgp_core_050;
  assign cgp_core_070 = input_f[0] & input_d[1];
  assign cgp_core_071 = ~cgp_core_046;
  assign cgp_core_072 = cgp_core_023 & cgp_core_071;
  assign cgp_core_073 = input_g[0] & input_b[1];
  assign cgp_core_074 = ~(cgp_core_023 ^ input_d[1]);
  assign cgp_core_075 = ~(cgp_core_074 | cgp_core_070);
  assign cgp_core_077 = cgp_core_059 ^ cgp_core_075;
  assign cgp_core_078 = cgp_core_063 | cgp_core_077;

  assign cgp_out[0] = 1'b0;
endmodule