module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, input [1:0] input_h, output [0:0] cgp_out);
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046_not;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052_not;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076_not;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_081_not;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_090;
  wire cgp_core_091;

  assign cgp_core_018 = input_f[0] ^ input_h[0];
  assign cgp_core_019 = ~(input_g[1] & input_a[0]);
  assign cgp_core_020 = ~input_h[0];
  assign cgp_core_021 = ~input_b[1];
  assign cgp_core_023 = input_c[0] & cgp_core_019;
  assign cgp_core_024 = cgp_core_021 & input_a[1];
  assign cgp_core_026 = ~(input_c[1] | input_e[0]);
  assign cgp_core_027 = input_a[1] ^ input_b[1];
  assign cgp_core_028 = ~(input_a[1] & input_c[0]);
  assign cgp_core_029 = ~(input_f[0] ^ input_d[0]);
  assign cgp_core_032 = input_b[0] | input_d[1];
  assign cgp_core_034 = ~(input_a[1] | input_h[0]);
  assign cgp_core_035 = input_h[0] & input_b[1];
  assign cgp_core_038 = ~(input_g[1] & input_a[1]);
  assign cgp_core_041 = ~(input_d[0] & cgp_core_034);
  assign cgp_core_042 = input_e[1] & cgp_core_034;
  assign cgp_core_043 = ~input_d[1];
  assign cgp_core_044 = input_d[1] & input_d[0];
  assign cgp_core_045 = ~(cgp_core_043 | input_e[1]);
  assign cgp_core_046_not = ~input_h[0];
  assign cgp_core_048 = input_b[1] ^ input_e[0];
  assign cgp_core_049 = input_a[0] & input_h[0];
  assign cgp_core_050 = ~input_g[1];
  assign cgp_core_052_not = ~input_e[1];
  assign cgp_core_054 = input_e[1] ^ input_c[0];
  assign cgp_core_055 = ~(input_c[0] & input_h[0]);
  assign cgp_core_057 = ~(input_c[1] & input_b[0]);
  assign cgp_core_061 = input_a[1] | input_d[0];
  assign cgp_core_063 = input_g[0] & input_f[0];
  assign cgp_core_065 = ~(input_b[1] & input_h[1]);
  assign cgp_core_066 = cgp_core_063 | cgp_core_065;
  assign cgp_core_067 = ~(input_e[0] & input_c[1]);
  assign cgp_core_069 = input_g[0] & input_b[0];
  assign cgp_core_070 = input_e[1] | input_f[1];
  assign cgp_core_071 = input_e[1] ^ input_c[0];
  assign cgp_core_073 = ~(cgp_core_070 & input_h[0]);
  assign cgp_core_074 = cgp_core_066 ^ cgp_core_066;
  assign cgp_core_076_not = ~input_d[0];
  assign cgp_core_078 = ~input_c[0];
  assign cgp_core_079 = input_b[0] & input_b[1];
  assign cgp_core_081_not = ~input_c[1];
  assign cgp_core_083 = ~input_b[1];
  assign cgp_core_085 = ~(input_e[1] ^ input_a[1]);
  assign cgp_core_086 = input_a[1] ^ input_b[0];
  assign cgp_core_090 = input_h[1] | input_c[0];
  assign cgp_core_091 = cgp_core_050 & cgp_core_067;

  assign cgp_out[0] = 1'b1;
endmodule