module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_038_not;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043_not;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_056_not;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_061_not;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_093_not;
  wire cgp_core_098;
  wire cgp_core_099;

  assign cgp_core_020 = input_e[0] & input_b[0];
  assign cgp_core_021 = ~(input_b[2] ^ input_a[0]);
  assign cgp_core_022 = ~(input_c[1] ^ input_b[2]);
  assign cgp_core_024 = input_e[1] | input_e[2];
  assign cgp_core_026 = input_c[2] & input_c[1];
  assign cgp_core_027 = input_c[2] | input_e[2];
  assign cgp_core_028 = input_c[2] & input_e[2];
  assign cgp_core_030 = cgp_core_027 & input_e[1];
  assign cgp_core_031 = cgp_core_028 | cgp_core_030;
  assign cgp_core_032 = ~(input_f[2] & input_c[1]);
  assign cgp_core_033 = input_c[0] | input_e[1];
  assign cgp_core_038_not = ~input_c[0];
  assign cgp_core_039 = input_d[0] & input_c[0];
  assign cgp_core_041 = ~input_f[2];
  assign cgp_core_043_not = ~input_e[2];
  assign cgp_core_045 = cgp_core_031 & input_a[2];
  assign cgp_core_046 = input_f[1] & input_b[2];
  assign cgp_core_047 = input_e[2] & input_b[2];
  assign cgp_core_049 = ~input_d[1];
  assign cgp_core_051 = ~(input_c[0] & input_b[1]);
  assign cgp_core_056_not = ~input_a[2];
  assign cgp_core_057 = input_c[0] & input_b[1];
  assign cgp_core_059 = input_e[1] & input_f[2];
  assign cgp_core_061_not = ~input_a[2];
  assign cgp_core_063 = ~(input_e[0] | input_a[1]);
  assign cgp_core_065 = input_f[0] | input_f[2];
  assign cgp_core_067 = ~(input_d[2] ^ input_f[1]);
  assign cgp_core_068 = input_d[0] | input_b[2];
  assign cgp_core_069_not = ~input_d[1];
  assign cgp_core_070 = input_d[2] & input_f[2];
  assign cgp_core_071 = ~input_f[0];
  assign cgp_core_072 = ~(input_e[0] & input_a[2]);
  assign cgp_core_074 = ~(input_e[1] | input_a[0]);
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = cgp_core_031 & cgp_core_075;
  assign cgp_core_078 = ~(input_b[2] | input_d[2]);
  assign cgp_core_080 = ~(input_c[1] ^ input_a[2]);
  assign cgp_core_082 = input_a[2] & cgp_core_078;
  assign cgp_core_083 = ~(input_b[2] ^ input_b[2]);
  assign cgp_core_084 = input_a[2] & input_d[1];
  assign cgp_core_085 = input_b[0] ^ input_c[1];
  assign cgp_core_086 = ~(input_b[1] ^ input_f[1]);
  assign cgp_core_087 = input_e[0] | input_f[0];
  assign cgp_core_088 = input_d[1] | input_f[1];
  assign cgp_core_090 = input_b[0] & input_c[2];
  assign cgp_core_093_not = ~input_b[0];
  assign cgp_core_098 = cgp_core_076 | cgp_core_045;
  assign cgp_core_099 = cgp_core_082 | cgp_core_098;

  assign cgp_out[0] = cgp_core_099;
endmodule