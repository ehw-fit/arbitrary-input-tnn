module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039_not;
  wire cgp_core_040_not;
  wire cgp_core_041;
  wire cgp_core_042_not;
  wire cgp_core_043;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = ~input_a[1];
  assign cgp_core_018 = input_a[2] & input_e[2];
  assign cgp_core_020 = ~input_a[2];
  assign cgp_core_022 = input_b[1] | input_a[0];
  assign cgp_core_024 = ~(input_b[0] & input_b[0]);
  assign cgp_core_025 = ~input_b[0];
  assign cgp_core_026 = input_c[1] | input_c[2];
  assign cgp_core_027 = input_b[1] | input_a[2];
  assign cgp_core_028 = input_d[0] ^ input_d[2];
  assign cgp_core_031 = input_b[1] & input_d[0];
  assign cgp_core_032 = input_b[1] & input_d[1];
  assign cgp_core_033 = ~(input_a[0] & input_b[1]);
  assign cgp_core_036 = input_a[1] & input_e[1];
  assign cgp_core_037 = input_b[1] | input_a[0];
  assign cgp_core_038 = input_b[2] | cgp_core_032;
  assign cgp_core_039_not = ~input_a[1];
  assign cgp_core_040_not = ~input_b[2];
  assign cgp_core_041 = ~(input_c[2] | input_a[0]);
  assign cgp_core_042_not = ~input_d[0];
  assign cgp_core_043 = input_e[0] ^ input_c[2];
  assign cgp_core_045 = input_d[1] ^ input_e[2];
  assign cgp_core_047 = ~input_c[1];
  assign cgp_core_048 = cgp_core_026 | cgp_core_038;
  assign cgp_core_049 = ~(input_b[2] | input_c[1]);
  assign cgp_core_050 = cgp_core_048 | input_d[2];
  assign cgp_core_051 = input_c[0] & input_b[0];
  assign cgp_core_054 = ~input_d[1];
  assign cgp_core_056 = input_c[1] ^ input_b[1];
  assign cgp_core_058 = input_a[0] & input_d[1];
  assign cgp_core_059 = input_d[0] ^ input_b[0];
  assign cgp_core_060 = ~input_e[0];
  assign cgp_core_061 = ~input_e[2];
  assign cgp_core_063 = ~cgp_core_050;
  assign cgp_core_064 = input_a[2] & cgp_core_063;
  assign cgp_core_065 = cgp_core_064 & cgp_core_061;
  assign cgp_core_068 = ~(input_d[2] ^ input_b[1]);
  assign cgp_core_069 = ~(input_d[2] | input_a[2]);
  assign cgp_core_071 = input_b[0] ^ input_a[1];
  assign cgp_core_072 = ~(input_e[2] ^ input_e[2]);
  assign cgp_core_073 = ~(input_a[2] | input_e[1]);
  assign cgp_core_074 = ~(input_c[1] & input_a[0]);
  assign cgp_core_076 = input_d[2] | input_d[2];
  assign cgp_core_077 = input_b[2] & input_d[2];
  assign cgp_core_078 = input_b[0] | input_c[2];
  assign cgp_core_079 = ~(input_e[2] & input_c[0]);

  assign cgp_out[0] = cgp_core_065;
endmodule