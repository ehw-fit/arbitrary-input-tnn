module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_029;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_036;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051_not;
  wire cgp_core_052;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;

  assign cgp_core_014 = input_a[0] ^ input_c[0];
  assign cgp_core_015 = input_f[0] & input_b[1];
  assign cgp_core_016 = input_a[1] ^ input_d[1];
  assign cgp_core_017 = input_d[1] & input_f[0];
  assign cgp_core_018 = input_c[1] ^ cgp_core_015;
  assign cgp_core_021 = input_e[0] & input_d[1];
  assign cgp_core_022 = input_e[0] & input_b[1];
  assign cgp_core_023 = input_a[1] & input_e[1];
  assign cgp_core_024 = ~input_e[0];
  assign cgp_core_026 = input_e[0] ^ cgp_core_022;
  assign cgp_core_027 = cgp_core_024 | cgp_core_026;
  assign cgp_core_028_not = ~input_a[0];
  assign cgp_core_029 = ~input_d[0];
  assign cgp_core_032 = ~(input_d[0] | cgp_core_029);
  assign cgp_core_033 = ~input_d[0];
  assign cgp_core_036 = input_f[0] & input_c[1];
  assign cgp_core_040 = input_b[0] | input_d[0];
  assign cgp_core_041 = input_c[0] ^ input_e[0];
  assign cgp_core_046 = input_b[0] | input_b[0];
  assign cgp_core_049 = ~(cgp_core_036 ^ input_b[0]);
  assign cgp_core_050 = input_d[1] ^ input_c[0];
  assign cgp_core_051_not = ~cgp_core_050;
  assign cgp_core_052 = input_d[0] | input_d[0];
  assign cgp_core_056 = input_a[1] ^ input_f[1];
  assign cgp_core_058 = ~input_b[0];
  assign cgp_core_059 = ~(input_a[1] | cgp_core_058);
  assign cgp_core_060 = cgp_core_059 | input_a[0];
  assign cgp_core_063 = input_e[1] & input_f[1];
  assign cgp_core_065 = ~(input_b[1] ^ input_b[0]);
  assign cgp_core_066 = ~(input_a[1] ^ input_e[1]);
  assign cgp_core_067 = input_f[1] & input_b[0];
  assign cgp_core_068 = ~(cgp_core_060 & input_f[1]);
  assign cgp_core_069 = input_e[1] | input_b[0];
  assign cgp_core_070 = input_e[1] | input_c[1];

  assign cgp_out[0] = 1'b1;
endmodule