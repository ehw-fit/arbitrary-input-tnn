module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_021;
  wire cgp_core_023_not;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_028;
  wire cgp_core_030_not;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_039_not;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;

  assign cgp_core_011 = input_b[2] & input_c[0];
  assign cgp_core_012 = ~(input_b[2] ^ input_c[0]);
  assign cgp_core_013 = ~(input_c[1] | input_a[0]);
  assign cgp_core_014 = ~input_b[0];
  assign cgp_core_016 = input_c[1] ^ input_b[0];
  assign cgp_core_017 = input_a[1] | input_c[0];
  assign cgp_core_021 = input_c[2] & input_a[0];
  assign cgp_core_023_not = ~input_b[0];
  assign cgp_core_024 = ~(input_a[0] ^ input_c[2]);
  assign cgp_core_025 = input_b[1] & input_a[1];
  assign cgp_core_028 = ~(input_b[2] | input_a[2]);
  assign cgp_core_030_not = ~input_c[2];
  assign cgp_core_031 = input_a[1] & input_c[2];
  assign cgp_core_032 = ~input_b[1];
  assign cgp_core_033_not = ~input_c[1];
  assign cgp_core_034 = input_a[0] & input_c[0];
  assign cgp_core_036 = ~(input_b[2] | input_b[1]);
  assign cgp_core_038 = input_a[2] & input_b[0];
  assign cgp_core_039_not = ~input_a[1];
  assign cgp_core_040 = input_b[2] | input_c[2];
  assign cgp_core_041 = cgp_core_025 | input_b[2];
  assign cgp_core_042 = input_a[2] | cgp_core_041;

  assign cgp_out[0] = cgp_core_042;
endmodule