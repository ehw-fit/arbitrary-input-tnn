module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_015;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_038;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044_not;
  wire cgp_core_045_not;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_070;

  assign cgp_core_015 = input_e[1] & input_c[0];
  assign cgp_core_017 = ~(input_c[1] | input_c[0]);
  assign cgp_core_018 = ~input_c[0];
  assign cgp_core_019 = input_a[1] & cgp_core_015;
  assign cgp_core_020 = input_f[1] | cgp_core_019;
  assign cgp_core_021 = input_f[0] ^ input_f[0];
  assign cgp_core_022 = input_e[0] & input_f[0];
  assign cgp_core_023 = input_c[0] ^ input_f[1];
  assign cgp_core_024 = input_f[1] & input_c[1];
  assign cgp_core_025 = cgp_core_023 ^ cgp_core_022;
  assign cgp_core_026 = cgp_core_023 & cgp_core_022;
  assign cgp_core_028 = ~(input_e[1] & input_e[0]);
  assign cgp_core_029 = input_d[1] & cgp_core_021;
  assign cgp_core_030 = input_d[1] & input_c[1];
  assign cgp_core_031 = input_b[1] & cgp_core_025;
  assign cgp_core_032 = input_a[0] ^ cgp_core_029;
  assign cgp_core_034 = ~(cgp_core_031 ^ input_f[0]);
  assign cgp_core_036 = input_f[1] & cgp_core_034;
  assign cgp_core_038 = ~(input_c[0] ^ input_f[0]);
  assign cgp_core_040 = input_c[1] & input_a[0];
  assign cgp_core_042 = ~input_b[0];
  assign cgp_core_043 = cgp_core_040 | input_e[0];
  assign cgp_core_044_not = ~cgp_core_020;
  assign cgp_core_045_not = ~cgp_core_020;
  assign cgp_core_047 = input_a[0] & input_c[1];
  assign cgp_core_048 = cgp_core_045_not | cgp_core_047;
  assign cgp_core_049 = cgp_core_036 ^ cgp_core_048;
  assign cgp_core_051 = ~(input_e[0] | input_c[1]);
  assign cgp_core_052 = cgp_core_049 & cgp_core_051;
  assign cgp_core_053 = input_c[0] & cgp_core_049;
  assign cgp_core_057 = input_c[0] | cgp_core_053;
  assign cgp_core_058 = ~input_b[1];
  assign cgp_core_061 = input_d[1] & input_c[0];
  assign cgp_core_062 = input_c[1] ^ input_b[1];
  assign cgp_core_066 = ~(input_f[0] ^ input_f[1]);
  assign cgp_core_067 = input_a[0] | input_e[1];
  assign cgp_core_070 = input_c[1] | cgp_core_067;

  assign cgp_out[0] = 1'b1;
endmodule