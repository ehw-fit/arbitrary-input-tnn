module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_016_not;
  wire cgp_core_017_not;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024_not;
  wire cgp_core_027_not;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035_not;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_055_not;
  wire cgp_core_056_not;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078_not;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_087_not;
  wire cgp_core_090;

  assign cgp_core_016_not = ~input_a[2];
  assign cgp_core_017_not = ~input_a[5];
  assign cgp_core_019 = input_a[9] & input_a[8];
  assign cgp_core_020 = input_a[9] | input_a[6];
  assign cgp_core_021 = ~input_a[12];
  assign cgp_core_022 = ~(input_a[12] ^ input_a[7]);
  assign cgp_core_024_not = ~input_a[10];
  assign cgp_core_027_not = ~input_a[9];
  assign cgp_core_028 = input_a[12] | input_a[5];
  assign cgp_core_029 = input_a[10] ^ input_a[13];
  assign cgp_core_030 = input_a[0] ^ input_a[11];
  assign cgp_core_031 = ~(input_a[4] & input_a[10]);
  assign cgp_core_032 = ~input_a[2];
  assign cgp_core_033 = ~(input_a[12] ^ input_a[7]);
  assign cgp_core_034 = input_a[1] | input_a[5];
  assign cgp_core_035_not = ~input_a[12];
  assign cgp_core_037 = input_a[10] | input_a[7];
  assign cgp_core_040 = input_a[11] ^ input_a[3];
  assign cgp_core_041 = input_a[11] ^ input_a[8];
  assign cgp_core_042 = ~(input_a[8] & input_a[5]);
  assign cgp_core_044 = ~(input_a[0] ^ input_a[10]);
  assign cgp_core_047 = ~(input_a[10] & input_a[10]);
  assign cgp_core_048 = ~(input_a[2] ^ input_a[8]);
  assign cgp_core_049 = input_a[9] ^ input_a[6];
  assign cgp_core_050 = ~(input_a[9] & input_a[13]);
  assign cgp_core_051 = ~(input_a[1] & input_a[1]);
  assign cgp_core_052 = ~(input_a[3] ^ input_a[7]);
  assign cgp_core_055_not = ~input_a[9];
  assign cgp_core_056_not = ~input_a[2];
  assign cgp_core_057 = ~input_a[5];
  assign cgp_core_058 = ~input_a[13];
  assign cgp_core_059 = input_a[12] | input_a[0];
  assign cgp_core_065 = ~(input_a[12] ^ input_a[3]);
  assign cgp_core_066 = input_a[12] & input_a[0];
  assign cgp_core_068 = ~(input_a[2] & input_a[10]);
  assign cgp_core_069 = input_a[7] | input_a[11];
  assign cgp_core_070 = ~input_a[4];
  assign cgp_core_072 = ~input_a[10];
  assign cgp_core_074 = input_a[9] & input_a[12];
  assign cgp_core_075 = ~(input_a[4] | input_a[12]);
  assign cgp_core_077 = input_a[8] ^ input_a[6];
  assign cgp_core_078_not = ~input_a[10];
  assign cgp_core_080 = ~input_a[1];
  assign cgp_core_082 = ~(input_a[10] & input_a[5]);
  assign cgp_core_083 = input_a[2] ^ input_a[13];
  assign cgp_core_085 = ~(input_a[1] | input_a[3]);
  assign cgp_core_087_not = ~input_a[1];
  assign cgp_core_090 = ~(input_a[0] | input_a[12]);

  assign cgp_out[0] = input_a[2];
  assign cgp_out[1] = 1'b1;
  assign cgp_out[2] = 1'b1;
  assign cgp_out[3] = 1'b0;
endmodule