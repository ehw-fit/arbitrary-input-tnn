module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048_not;
  wire cgp_core_050_not;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_066_not;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = ~(input_d[0] | input_b[0]);
  assign cgp_core_018 = ~input_c[2];
  assign cgp_core_019 = ~(input_b[1] | input_e[2]);
  assign cgp_core_021 = cgp_core_019 ^ input_a[2];
  assign cgp_core_022 = ~(input_d[0] ^ input_a[1]);
  assign cgp_core_029 = ~(input_a[1] | input_c[1]);
  assign cgp_core_030 = input_a[2] & input_b[0];
  assign cgp_core_032 = ~(input_d[1] & input_e[1]);
  assign cgp_core_035 = ~input_a[0];
  assign cgp_core_036 = input_d[1] ^ input_e[1];
  assign cgp_core_037 = ~input_c[1];
  assign cgp_core_040 = input_a[2] & input_d[1];
  assign cgp_core_041 = ~(input_c[2] | input_d[1]);
  assign cgp_core_042 = ~(cgp_core_017 & input_a[1]);
  assign cgp_core_045 = ~(input_d[0] & input_e[0]);
  assign cgp_core_046 = input_c[2] & input_e[1];
  assign cgp_core_048_not = ~input_b[0];
  assign cgp_core_050_not = ~input_e[1];
  assign cgp_core_051 = ~(input_e[1] ^ input_b[0]);
  assign cgp_core_053 = input_a[2] ^ input_d[0];
  assign cgp_core_054 = ~(input_a[2] ^ input_b[0]);
  assign cgp_core_055 = ~(input_e[1] & input_e[1]);
  assign cgp_core_057 = ~input_c[1];
  assign cgp_core_059 = input_c[0] | input_b[1];
  assign cgp_core_061 = ~(input_e[0] & input_b[1]);
  assign cgp_core_066_not = ~input_d[1];
  assign cgp_core_067 = ~(input_b[2] & input_e[0]);
  assign cgp_core_068 = input_c[0] ^ cgp_core_045;
  assign cgp_core_069 = ~(input_c[0] & input_a[0]);
  assign cgp_core_070 = input_a[1] ^ input_b[0];
  assign cgp_core_071 = ~(input_a[0] | input_a[1]);
  assign cgp_core_074 = ~(input_b[2] & input_b[1]);
  assign cgp_core_075 = input_d[0] & input_d[1];
  assign cgp_core_076 = ~(input_d[2] & input_c[1]);
  assign cgp_core_077 = input_a[0] & input_a[2];
  assign cgp_core_078 = ~(input_a[2] | input_b[1]);
  assign cgp_core_079 = ~input_d[0];

  assign cgp_out[0] = 1'b0;
endmodule