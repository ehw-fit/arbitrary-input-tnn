module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015_not;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_047;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_058;

  assign cgp_core_014 = ~input_d[2];
  assign cgp_core_015_not = ~input_d[0];
  assign cgp_core_016 = ~(input_a[0] & input_b[0]);
  assign cgp_core_017 = input_a[1] & input_b[1];
  assign cgp_core_018 = input_c[0] | input_a[2];
  assign cgp_core_021 = input_a[2] | input_b[2];
  assign cgp_core_022 = input_a[2] & input_b[2];
  assign cgp_core_023 = input_d[0] | input_b[1];
  assign cgp_core_024 = cgp_core_021 & cgp_core_017;
  assign cgp_core_025 = cgp_core_022 | cgp_core_024;
  assign cgp_core_026 = ~(input_b[2] ^ input_d[2]);
  assign cgp_core_027 = input_d[0] & input_a[0];
  assign cgp_core_028 = input_d[2] & input_d[2];
  assign cgp_core_029 = input_a[2] ^ input_b[0];
  assign cgp_core_030 = ~(input_b[2] | input_d[0]);
  assign cgp_core_031 = input_a[2] ^ input_c[0];
  assign cgp_core_033 = input_c[2] | input_d[2];
  assign cgp_core_034 = ~(input_c[0] & input_b[1]);
  assign cgp_core_036 = ~(input_c[0] & input_b[1]);
  assign cgp_core_041 = ~cgp_core_033;
  assign cgp_core_044 = input_b[0] ^ input_d[1];
  assign cgp_core_047 = ~input_d[1];
  assign cgp_core_049_not = ~input_b[0];
  assign cgp_core_050 = ~(input_d[1] & input_d[0]);
  assign cgp_core_058 = cgp_core_041 | cgp_core_025;

  assign cgp_out[0] = cgp_core_058;
endmodule