module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, input [2:0] input_f, output [0:0] cgp_out);
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023_not;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_081;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_096;
  wire cgp_core_098;

  assign cgp_core_021 = ~(input_c[1] & input_c[2]);
  assign cgp_core_022 = ~(input_a[0] ^ input_d[1]);
  assign cgp_core_023_not = ~input_d[0];
  assign cgp_core_026 = input_c[0] | input_f[0];
  assign cgp_core_028 = ~(input_a[1] ^ input_f[2]);
  assign cgp_core_029 = input_d[2] & input_a[0];
  assign cgp_core_030 = ~(input_a[2] ^ input_b[2]);
  assign cgp_core_031 = input_e[2] | input_c[2];
  assign cgp_core_032 = ~input_c[2];
  assign cgp_core_033 = ~input_a[0];
  assign cgp_core_034 = ~input_e[1];
  assign cgp_core_036 = ~(input_f[0] & input_a[2]);
  assign cgp_core_037 = ~(input_a[0] | input_e[2]);
  assign cgp_core_038 = ~(input_d[2] & input_c[1]);
  assign cgp_core_039 = input_a[1] | input_e[1];
  assign cgp_core_043 = input_a[2] | cgp_core_039;
  assign cgp_core_044 = ~(input_b[0] | input_c[1]);
  assign cgp_core_045 = cgp_core_031 & cgp_core_043;
  assign cgp_core_046 = input_b[0] | input_c[1];
  assign cgp_core_050 = input_c[1] | input_b[2];
  assign cgp_core_051 = ~input_e[1];
  assign cgp_core_053 = ~(input_c[0] | input_a[2]);
  assign cgp_core_054 = input_d[2] & input_f[2];
  assign cgp_core_056 = ~input_d[2];
  assign cgp_core_058 = ~input_f[2];
  assign cgp_core_061 = ~(input_f[2] & input_f[1]);
  assign cgp_core_063 = input_c[0] ^ input_d[0];
  assign cgp_core_064 = ~input_e[2];
  assign cgp_core_065 = ~input_e[1];
  assign cgp_core_066 = ~(input_f[2] & input_b[2]);
  assign cgp_core_067 = ~(input_e[2] | input_a[0]);
  assign cgp_core_068 = ~(input_c[1] ^ input_c[1]);
  assign cgp_core_070 = input_b[2] | input_f[2];
  assign cgp_core_071 = cgp_core_054 & input_b[2];
  assign cgp_core_072 = ~cgp_core_071;
  assign cgp_core_073 = cgp_core_045 & cgp_core_072;
  assign cgp_core_075 = ~cgp_core_070;
  assign cgp_core_076 = input_c[1] & cgp_core_075;
  assign cgp_core_078 = input_a[1] & input_f[0];
  assign cgp_core_081 = ~input_e[1];
  assign cgp_core_084 = input_d[2] ^ input_f[0];
  assign cgp_core_085 = ~(input_a[2] ^ input_b[2]);
  assign cgp_core_086 = ~(input_f[1] ^ input_c[0]);
  assign cgp_core_088 = ~input_f[0];
  assign cgp_core_092 = ~input_d[0];
  assign cgp_core_093 = ~input_c[2];
  assign cgp_core_096 = ~input_a[2];
  assign cgp_core_098 = cgp_core_076 | cgp_core_073;

  assign cgp_out[0] = cgp_core_098;
endmodule