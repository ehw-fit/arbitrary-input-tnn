module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, input [1:0] input_g, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_034;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_046;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052_not;
  wire cgp_core_054;
  wire cgp_core_057_not;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065_not;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;

  assign cgp_core_017 = input_c[0] & input_e[0];
  assign cgp_core_018 = input_b[0] ^ input_a[1];
  assign cgp_core_019 = input_c[1] & input_d[0];
  assign cgp_core_022 = cgp_core_019 & input_e[0];
  assign cgp_core_024 = ~(input_a[0] & input_g[0]);
  assign cgp_core_025 = ~(input_d[0] & input_c[1]);
  assign cgp_core_026 = ~(input_a[1] | input_f[0]);
  assign cgp_core_028 = ~(input_d[1] ^ cgp_core_024);
  assign cgp_core_029 = ~input_g[1];
  assign cgp_core_030 = input_g[0] | input_d[0];
  assign cgp_core_031 = ~(cgp_core_022 & input_g[1]);
  assign cgp_core_034 = input_f[0] & input_d[1];
  assign cgp_core_039 = input_f[0] ^ input_g[1];
  assign cgp_core_041 = ~input_a[0];
  assign cgp_core_043 = cgp_core_041 ^ input_d[1];
  assign cgp_core_046 = input_e[1] & input_c[0];
  assign cgp_core_049 = ~(input_f[0] ^ input_c[0]);
  assign cgp_core_050 = ~input_c[0];
  assign cgp_core_052_not = ~cgp_core_049;
  assign cgp_core_054 = input_a[0] | input_e[0];
  assign cgp_core_057_not = ~input_g[1];
  assign cgp_core_058 = input_g[0] | input_a[1];
  assign cgp_core_060 = input_d[1] & cgp_core_057_not;
  assign cgp_core_062 = ~(input_a[0] | input_d[0]);
  assign cgp_core_063 = ~(input_f[1] & input_e[0]);
  assign cgp_core_065_not = ~input_b[1];
  assign cgp_core_068 = ~(input_c[1] ^ input_g[0]);
  assign cgp_core_069 = ~(input_c[0] ^ input_g[0]);
  assign cgp_core_073 = input_e[0] & input_c[1];
  assign cgp_core_074 = input_f[0] ^ cgp_core_046;
  assign cgp_core_076 = cgp_core_073 & input_a[0];
  assign cgp_core_078 = input_g[1] | input_d[1];
  assign cgp_core_079 = ~(input_f[0] & input_d[0]);

  assign cgp_out[0] = input_d[0];
endmodule