module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, output [0:0] cgp_out);
  wire cgp_core_011;
  wire cgp_core_012;
  wire cgp_core_013;
  wire cgp_core_014;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_027;
  wire cgp_core_029_not;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_042;

  assign cgp_core_011 = ~input_c[1];
  assign cgp_core_012 = ~(input_b[0] ^ input_b[0]);
  assign cgp_core_013 = input_b[0] ^ input_a[1];
  assign cgp_core_014 = ~(input_c[0] | input_b[2]);
  assign cgp_core_017 = input_c[1] ^ input_c[2];
  assign cgp_core_018 = input_b[2] | input_b[1];
  assign cgp_core_019 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_020 = input_b[2] | input_b[1];
  assign cgp_core_021 = input_b[2] & input_b[1];
  assign cgp_core_022 = input_a[2] | cgp_core_021;
  assign cgp_core_024 = ~input_c[2];
  assign cgp_core_025 = cgp_core_020 & cgp_core_024;
  assign cgp_core_027 = ~(input_b[2] ^ input_c[2]);
  assign cgp_core_029_not = ~input_c[2];
  assign cgp_core_031 = input_a[1] & cgp_core_027;
  assign cgp_core_033 = ~(input_a[2] & input_a[1]);
  assign cgp_core_034 = ~(input_b[2] & input_b[0]);
  assign cgp_core_035 = input_c[2] ^ input_b[1];
  assign cgp_core_037 = ~input_b[0];
  assign cgp_core_038 = input_c[0] ^ input_b[2];
  assign cgp_core_041 = cgp_core_025 | cgp_core_022;
  assign cgp_core_042 = cgp_core_031 | cgp_core_041;

  assign cgp_out[0] = cgp_core_042;
endmodule