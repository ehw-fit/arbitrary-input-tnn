module cgp(input [11:0] input_a, output [3:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_023;
  wire cgp_core_027;
  wire cgp_core_029;
  wire cgp_core_034_not;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_042;
  wire cgp_core_045;
  wire cgp_core_049;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_078;

  assign cgp_core_014 = ~(input_a[11] | input_a[1]);
  assign cgp_core_015 = input_a[2] ^ input_a[3];
  assign cgp_core_016 = ~input_a[4];
  assign cgp_core_019 = ~(input_a[9] ^ input_a[5]);
  assign cgp_core_020 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_021 = input_a[9] & input_a[7];
  assign cgp_core_022 = ~input_a[2];
  assign cgp_core_023 = ~(input_a[9] ^ input_a[7]);
  assign cgp_core_027 = ~(input_a[7] ^ input_a[8]);
  assign cgp_core_029 = input_a[3] & input_a[11];
  assign cgp_core_034_not = ~input_a[9];
  assign cgp_core_035 = ~(input_a[11] & input_a[0]);
  assign cgp_core_037 = ~(input_a[3] & input_a[1]);
  assign cgp_core_038 = ~input_a[6];
  assign cgp_core_039 = input_a[6] ^ input_a[5];
  assign cgp_core_042 = ~(input_a[8] | input_a[7]);
  assign cgp_core_045 = ~input_a[10];
  assign cgp_core_049 = input_a[8] & input_a[11];
  assign cgp_core_055 = ~(input_a[3] & input_a[6]);
  assign cgp_core_057 = input_a[6] ^ input_a[1];
  assign cgp_core_062 = input_a[6] & input_a[4];
  assign cgp_core_064 = ~input_a[3];
  assign cgp_core_065 = ~(input_a[7] ^ input_a[2]);
  assign cgp_core_067 = input_a[3] ^ input_a[0];
  assign cgp_core_068 = input_a[9] | input_a[4];
  assign cgp_core_072 = ~input_a[2];
  assign cgp_core_073 = input_a[7] | input_a[1];
  assign cgp_core_074 = ~(input_a[0] & input_a[3]);
  assign cgp_core_078 = ~(input_a[7] & input_a[1]);

  assign cgp_out[0] = 1'b0;
  assign cgp_out[1] = 1'b0;
  assign cgp_out[2] = 1'b0;
  assign cgp_out[3] = 1'b1;
endmodule