module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033_not;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064_not;
  wire cgp_core_065;
  wire cgp_core_066_not;
  wire cgp_core_070;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017 = ~(input_a[0] ^ input_a[1]);
  assign cgp_core_019 = ~(input_d[2] ^ input_c[1]);
  assign cgp_core_020 = input_b[2] | input_e[1];
  assign cgp_core_021 = ~(input_d[0] | input_d[1]);
  assign cgp_core_024 = input_e[1] ^ input_b[1];
  assign cgp_core_025 = ~(input_c[0] & input_d[0]);
  assign cgp_core_026 = input_a[0] | input_a[0];
  assign cgp_core_027 = input_c[1] | input_e[0];
  assign cgp_core_028 = input_a[2] ^ input_e[1];
  assign cgp_core_031 = ~(input_a[0] & input_e[1]);
  assign cgp_core_032 = ~input_e[2];
  assign cgp_core_033_not = ~input_e[2];
  assign cgp_core_034 = input_c[2] ^ input_b[1];
  assign cgp_core_035 = input_d[1] ^ input_d[1];
  assign cgp_core_038 = input_e[1] | input_c[0];
  assign cgp_core_039 = input_c[2] ^ input_e[2];
  assign cgp_core_040 = input_a[0] ^ input_e[2];
  assign cgp_core_043 = ~(input_a[1] | input_a[2]);
  assign cgp_core_044 = input_d[0] & input_e[1];
  assign cgp_core_048 = input_c[0] & input_a[0];
  assign cgp_core_049 = input_a[2] | input_c[1];
  assign cgp_core_051 = input_a[2] | input_c[1];
  assign cgp_core_052 = ~input_a[1];
  assign cgp_core_053 = ~(input_a[0] & input_b[2]);
  assign cgp_core_055 = input_b[2] & input_a[1];
  assign cgp_core_057 = ~(input_e[2] | input_b[1]);
  assign cgp_core_058 = ~(input_a[2] ^ input_d[1]);
  assign cgp_core_059 = ~(input_d[1] ^ input_e[0]);
  assign cgp_core_060 = ~input_a[2];
  assign cgp_core_061 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_063 = input_a[0] & input_a[2];
  assign cgp_core_064_not = ~input_d[2];
  assign cgp_core_065 = ~(input_e[2] | input_b[2]);
  assign cgp_core_066_not = ~input_a[2];
  assign cgp_core_070 = ~(input_d[1] & input_c[2]);
  assign cgp_core_073 = ~input_a[0];
  assign cgp_core_074 = input_d[2] | input_a[2];
  assign cgp_core_075 = input_c[2] | input_c[2];
  assign cgp_core_079 = input_b[2] | input_e[2];
  assign cgp_core_080 = input_c[2] | cgp_core_079;

  assign cgp_out[0] = cgp_core_080;
endmodule