module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_022_not;
  wire cgp_core_023;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_037;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_048;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_017 = input_a[1] ^ input_e[0];
  assign cgp_core_018 = input_c[2] & input_d[0];
  assign cgp_core_019 = ~(input_a[2] ^ input_c[0]);
  assign cgp_core_022_not = ~input_e[2];
  assign cgp_core_023 = input_c[0] ^ input_e[1];
  assign cgp_core_024 = ~(input_a[1] ^ input_b[2]);
  assign cgp_core_025 = input_e[0] & input_c[1];
  assign cgp_core_026 = input_b[0] & input_d[1];
  assign cgp_core_029 = input_e[0] | input_a[0];
  assign cgp_core_031 = ~(input_e[1] | input_b[1]);
  assign cgp_core_033 = input_d[0] ^ input_a[0];
  assign cgp_core_037 = ~(input_e[1] & input_a[0]);
  assign cgp_core_040 = input_e[1] | input_b[1];
  assign cgp_core_041 = input_d[1] & input_e[0];
  assign cgp_core_042 = ~(input_c[1] & input_e[1]);
  assign cgp_core_043 = ~(input_a[1] ^ input_e[1]);
  assign cgp_core_044 = ~(input_d[2] | input_d[0]);
  assign cgp_core_048 = input_e[2] ^ input_a[1];
  assign cgp_core_050 = input_a[1] ^ input_c[0];
  assign cgp_core_052 = input_b[0] ^ input_b[0];
  assign cgp_core_055 = ~(input_c[0] | input_b[2]);
  assign cgp_core_056 = ~(input_b[0] ^ input_b[0]);
  assign cgp_core_059 = ~(input_e[2] | input_b[0]);
  assign cgp_core_060 = ~(input_c[1] & input_e[1]);
  assign cgp_core_061 = input_d[0] & input_b[1];
  assign cgp_core_062 = ~(input_c[0] & input_d[0]);
  assign cgp_core_064 = input_a[2] & input_b[1];
  assign cgp_core_065 = ~(input_b[0] | input_c[2]);
  assign cgp_core_066 = ~(input_b[0] & input_d[2]);
  assign cgp_core_070 = ~(input_e[2] | input_b[1]);
  assign cgp_core_071 = ~(input_c[2] & input_b[0]);
  assign cgp_core_072 = ~input_c[0];
  assign cgp_core_074 = input_d[0] ^ input_c[0];
  assign cgp_core_075 = input_d[1] ^ input_a[2];
  assign cgp_core_076 = ~(input_a[1] ^ input_a[1]);
  assign cgp_core_078 = input_d[0] ^ input_a[0];
  assign cgp_core_079 = input_e[2] | input_c[2];
  assign cgp_core_080 = input_e[1] | cgp_core_079;

  assign cgp_out[0] = cgp_core_080;
endmodule