module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_018_not;
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034_not;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_041;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;

  assign cgp_core_018_not = ~input_a[0];
  assign cgp_core_019 = input_b[1] ^ input_c[1];
  assign cgp_core_020 = input_b[1] & input_c[1];
  assign cgp_core_024 = input_a[0] & input_d[0];
  assign cgp_core_025 = input_a[2] & input_e[2];
  assign cgp_core_026 = input_c[2] | cgp_core_020;
  assign cgp_core_027 = input_c[2] & input_c[1];
  assign cgp_core_028 = input_b[2] | cgp_core_027;
  assign cgp_core_029 = ~(input_d[0] | input_c[2]);
  assign cgp_core_030 = input_e[1] | input_d[1];
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_033 = input_d[1] | input_e[1];
  assign cgp_core_034_not = ~input_b[1];
  assign cgp_core_036 = input_a[0] & input_d[0];
  assign cgp_core_037 = ~(input_d[1] | input_b[2]);
  assign cgp_core_038 = input_e[2] | cgp_core_032;
  assign cgp_core_041 = input_a[1] ^ input_c[0];
  assign cgp_core_043 = cgp_core_019 ^ cgp_core_033;
  assign cgp_core_044 = cgp_core_019 & cgp_core_033;
  assign cgp_core_046 = ~input_c[2];
  assign cgp_core_048 = cgp_core_026 | cgp_core_038;
  assign cgp_core_049 = cgp_core_026 & input_e[2];
  assign cgp_core_050 = cgp_core_048 | cgp_core_044;
  assign cgp_core_051 = cgp_core_048 & cgp_core_044;
  assign cgp_core_052 = cgp_core_049 | cgp_core_051;
  assign cgp_core_053 = ~(input_a[2] | input_c[2]);
  assign cgp_core_055 = input_d[2] | cgp_core_052;
  assign cgp_core_059 = ~cgp_core_028;
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_062 = cgp_core_061 & cgp_core_059;
  assign cgp_core_063 = ~cgp_core_050;
  assign cgp_core_064 = input_a[2] & cgp_core_063;
  assign cgp_core_065 = cgp_core_064 & cgp_core_062;
  assign cgp_core_066 = ~(input_a[2] ^ cgp_core_050);
  assign cgp_core_067 = cgp_core_066 & cgp_core_062;
  assign cgp_core_068 = ~cgp_core_043;
  assign cgp_core_069 = input_a[1] & cgp_core_068;
  assign cgp_core_070 = cgp_core_069 & cgp_core_067;
  assign cgp_core_071 = ~(input_a[0] | input_b[1]);
  assign cgp_core_073 = ~input_e[2];
  assign cgp_core_074 = input_d[0] ^ input_a[2];
  assign cgp_core_076 = ~(input_c[2] | input_e[0]);
  assign cgp_core_077 = ~(input_e[2] | input_e[1]);
  assign cgp_core_078 = cgp_core_070 | cgp_core_065;
  assign cgp_core_079 = ~(input_b[0] & input_d[0]);
  assign cgp_core_080 = input_d[1] | input_a[2];

  assign cgp_out[0] = cgp_core_078;
endmodule