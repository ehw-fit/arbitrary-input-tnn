module cgp(input [1:0] input_a, input [1:0] input_b, input [1:0] input_c, input [1:0] input_d, input [1:0] input_e, input [1:0] input_f, output [0:0] cgp_out);
  wire cgp_core_014;
  wire cgp_core_015;
  wire cgp_core_016;
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_020;
  wire cgp_core_021;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_030_not;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_037_not;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_061;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_071;

  assign cgp_core_014 = input_d[1] ^ input_a[1];
  assign cgp_core_015 = input_f[0] & input_c[0];
  assign cgp_core_016 = ~(input_a[1] | input_b[0]);
  assign cgp_core_017 = input_e[1] & input_c[1];
  assign cgp_core_018 = cgp_core_016 | input_d[1];
  assign cgp_core_020 = ~(cgp_core_017 | input_f[1]);
  assign cgp_core_021 = ~(input_e[0] & input_f[0]);
  assign cgp_core_022 = ~(input_e[0] ^ input_f[0]);
  assign cgp_core_024 = input_f[0] & input_f[1];
  assign cgp_core_028 = ~(input_f[1] & cgp_core_021);
  assign cgp_core_029 = input_a[1] | cgp_core_021;
  assign cgp_core_030_not = ~input_c[1];
  assign cgp_core_031 = ~(input_d[1] | input_b[1]);
  assign cgp_core_032 = ~input_d[1];
  assign cgp_core_034 = ~input_e[1];
  assign cgp_core_037_not = ~input_d[1];
  assign cgp_core_039 = ~(input_c[0] | input_e[1]);
  assign cgp_core_041 = ~input_e[1];
  assign cgp_core_045 = ~(input_c[1] & cgp_core_024);
  assign cgp_core_047 = ~input_b[0];
  assign cgp_core_048 = cgp_core_045 | cgp_core_047;
  assign cgp_core_049 = input_e[0] | cgp_core_048;
  assign cgp_core_050 = input_a[1] & input_f[1];
  assign cgp_core_052 = ~(input_a[0] & input_b[0]);
  assign cgp_core_053 = ~input_c[0];
  assign cgp_core_058 = ~(input_f[1] | input_c[1]);
  assign cgp_core_059 = ~(input_f[0] | input_d[0]);
  assign cgp_core_061 = ~(input_f[0] ^ input_b[1]);
  assign cgp_core_064 = input_d[0] & input_f[0];
  assign cgp_core_065 = ~input_d[0];
  assign cgp_core_066 = ~input_c[1];
  assign cgp_core_071 = ~input_e[0];

  assign cgp_out[0] = 1'b1;
endmodule