module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_018;
  wire cgp_core_019;
  wire cgp_core_021;
  wire cgp_core_026;
  wire cgp_core_028;
  wire cgp_core_029;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_042;
  wire cgp_core_045_not;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_073;

  assign cgp_core_017 = input_b[0] ^ input_b[2];
  assign cgp_core_018 = input_c[1] & input_c[0];
  assign cgp_core_019 = input_b[0] ^ input_c[2];
  assign cgp_core_021 = cgp_core_019 ^ input_c[2];
  assign cgp_core_026 = ~input_b[2];
  assign cgp_core_028 = input_a[1] | input_b[2];
  assign cgp_core_029 = input_a[2] ^ input_e[0];
  assign cgp_core_031 = input_d[1] ^ input_e[1];
  assign cgp_core_032 = input_d[1] & input_e[1];
  assign cgp_core_034 = cgp_core_031 & input_d[0];
  assign cgp_core_035 = input_a[0] | input_b[1];
  assign cgp_core_037 = input_d[2] & input_e[2];
  assign cgp_core_038 = input_d[2] ^ input_c[1];
  assign cgp_core_039 = input_d[2] & cgp_core_035;
  assign cgp_core_040 = cgp_core_037 | input_a[2];
  assign cgp_core_042 = ~(cgp_core_017 | cgp_core_029);
  assign cgp_core_045_not = ~cgp_core_042;
  assign cgp_core_049 = cgp_core_026 & cgp_core_038;
  assign cgp_core_050 = cgp_core_026 ^ input_a[2];
  assign cgp_core_051 = ~cgp_core_026;
  assign cgp_core_052 = input_d[2] | cgp_core_051;
  assign cgp_core_053 = cgp_core_028 ^ cgp_core_040;
  assign cgp_core_054 = cgp_core_028 & cgp_core_040;
  assign cgp_core_055 = cgp_core_053 ^ cgp_core_052;
  assign cgp_core_056 = cgp_core_053 & cgp_core_052;
  assign cgp_core_057 = cgp_core_054 | cgp_core_056;
  assign cgp_core_058 = ~input_a[1];
  assign cgp_core_060 = ~cgp_core_055;
  assign cgp_core_061 = ~cgp_core_055;
  assign cgp_core_063 = ~cgp_core_050;
  assign cgp_core_064 = input_a[2] & input_b[0];
  assign cgp_core_066 = ~(input_a[2] ^ cgp_core_050);
  assign cgp_core_068 = cgp_core_045_not & cgp_core_045_not;
  assign cgp_core_069 = input_d[1] | input_e[1];
  assign cgp_core_071 = ~(input_a[1] ^ cgp_core_045_not);
  assign cgp_core_073 = ~input_e[2];

  assign cgp_out[0] = 1'b0;
endmodule