module cgp(input [13:0] input_a, output [3:0] cgp_out);
  wire cgp_core_017;
  wire cgp_core_021_not;
  wire cgp_core_023_not;
  wire cgp_core_026;
  wire cgp_core_031;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_068;
  wire cgp_core_069_not;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_083;
  wire cgp_core_086;
  wire cgp_core_087_not;
  wire cgp_core_088;
  wire cgp_core_089;

  assign cgp_core_017 = input_a[3] & input_a[9];
  assign cgp_core_021_not = ~input_a[4];
  assign cgp_core_023_not = ~input_a[7];
  assign cgp_core_026 = ~(input_a[12] ^ input_a[6]);
  assign cgp_core_031 = ~(input_a[1] & input_a[11]);
  assign cgp_core_033 = ~(input_a[5] | input_a[12]);
  assign cgp_core_035 = input_a[1] & input_a[6];
  assign cgp_core_036 = input_a[13] & input_a[4];
  assign cgp_core_037 = ~input_a[10];
  assign cgp_core_041 = input_a[8] & input_a[0];
  assign cgp_core_042 = ~(input_a[9] ^ input_a[8]);
  assign cgp_core_043 = ~(input_a[3] | input_a[9]);
  assign cgp_core_044 = input_a[12] ^ input_a[5];
  assign cgp_core_046 = ~(input_a[5] & input_a[10]);
  assign cgp_core_047 = input_a[1] ^ input_a[7];
  assign cgp_core_049 = ~(input_a[5] | input_a[13]);
  assign cgp_core_051 = ~input_a[1];
  assign cgp_core_052 = input_a[4] & input_a[8];
  assign cgp_core_053 = ~input_a[7];
  assign cgp_core_056 = ~input_a[5];
  assign cgp_core_057 = input_a[13] | input_a[12];
  assign cgp_core_060 = input_a[10] & input_a[10];
  assign cgp_core_063 = ~(input_a[7] | input_a[6]);
  assign cgp_core_064 = ~(input_a[7] ^ input_a[1]);
  assign cgp_core_065 = input_a[5] & input_a[12];
  assign cgp_core_068 = ~(input_a[13] | input_a[13]);
  assign cgp_core_069_not = ~input_a[1];
  assign cgp_core_070 = ~(input_a[3] & input_a[11]);
  assign cgp_core_071 = input_a[12] ^ input_a[9];
  assign cgp_core_072 = ~(input_a[9] ^ input_a[0]);
  assign cgp_core_074 = input_a[13] | input_a[2];
  assign cgp_core_075 = ~(input_a[6] & input_a[2]);
  assign cgp_core_078 = ~(input_a[0] ^ input_a[4]);
  assign cgp_core_079 = ~(input_a[8] ^ input_a[8]);
  assign cgp_core_080 = ~(input_a[13] ^ input_a[5]);
  assign cgp_core_081 = input_a[11] & input_a[7];
  assign cgp_core_083 = ~(input_a[9] | input_a[11]);
  assign cgp_core_086 = ~(input_a[4] | input_a[9]);
  assign cgp_core_087_not = ~input_a[13];
  assign cgp_core_088 = input_a[9] | input_a[13];
  assign cgp_core_089 = ~(input_a[12] ^ input_a[2]);

  assign cgp_out[0] = 1'b0;
  assign cgp_out[1] = 1'b1;
  assign cgp_out[2] = input_a[8];
  assign cgp_out[3] = input_a[2];
endmodule