module cgp(input [2:0] input_a, input [2:0] input_b, input [2:0] input_c, input [2:0] input_d, input [2:0] input_e, output [0:0] cgp_out);
  wire cgp_core_019;
  wire cgp_core_020;
  wire cgp_core_022;
  wire cgp_core_024;
  wire cgp_core_025;
  wire cgp_core_026;
  wire cgp_core_027;
  wire cgp_core_028_not;
  wire cgp_core_030;
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_039;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_049_not;
  wire cgp_core_050;
  wire cgp_core_053;
  wire cgp_core_056;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061_not;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;

  assign cgp_core_019 = ~input_e[0];
  assign cgp_core_020 = ~(input_e[1] & input_a[0]);
  assign cgp_core_022 = ~(cgp_core_019 & input_a[2]);
  assign cgp_core_024 = ~(input_c[2] & input_a[2]);
  assign cgp_core_025 = ~(input_c[2] & input_b[2]);
  assign cgp_core_026 = input_d[2] ^ input_e[0];
  assign cgp_core_027 = input_a[2] ^ input_c[0];
  assign cgp_core_028_not = ~input_a[0];
  assign cgp_core_030 = input_b[2] & input_e[1];
  assign cgp_core_031 = ~(input_b[1] & input_c[0]);
  assign cgp_core_032 = ~input_b[2];
  assign cgp_core_033 = ~(input_a[0] ^ input_e[2]);
  assign cgp_core_035 = ~input_a[1];
  assign cgp_core_037 = ~input_a[2];
  assign cgp_core_039 = input_a[2] | input_b[1];
  assign cgp_core_041 = input_d[0] | input_a[2];
  assign cgp_core_042 = ~input_a[0];
  assign cgp_core_043 = input_c[2] | input_b[1];
  assign cgp_core_044 = ~input_a[1];
  assign cgp_core_045 = input_c[2] ^ input_c[1];
  assign cgp_core_046 = ~input_e[0];
  assign cgp_core_047 = ~(input_b[0] ^ input_a[0]);
  assign cgp_core_049_not = ~input_d[0];
  assign cgp_core_050 = input_d[0] ^ input_d[2];
  assign cgp_core_053 = ~(input_e[1] ^ input_e[2]);
  assign cgp_core_056 = ~(input_c[0] & input_c[2]);
  assign cgp_core_058 = ~(input_a[2] | input_e[1]);
  assign cgp_core_060 = ~(input_b[1] & input_b[0]);
  assign cgp_core_061_not = ~input_b[0];
  assign cgp_core_067 = ~(input_c[1] ^ input_b[2]);
  assign cgp_core_068 = input_e[2] ^ input_e[0];
  assign cgp_core_069 = input_d[2] ^ input_c[1];
  assign cgp_core_076 = ~(input_d[2] ^ input_d[1]);
  assign cgp_core_077 = input_c[2] | input_d[0];
  assign cgp_core_079 = ~input_d[0];

  assign cgp_out[0] = 1'b1;
endmodule